magic
tech sky130A
timestamp 1620577694
<< nwell >>
rect 1010 1270 1215 1295
rect 990 1080 1215 1270
rect 1010 1055 1215 1080
rect 1200 395 1215 635
<< poly >>
rect 180 685 195 720
rect 180 670 400 685
rect 90 660 130 670
rect 90 640 100 660
rect 120 640 130 660
rect 90 630 130 640
rect 385 630 400 670
rect 1130 670 1170 680
rect 1130 650 1140 670
rect 1160 650 1170 670
rect 1130 640 1170 650
rect 1130 630 1145 640
<< polycont >>
rect 100 640 120 660
rect 1140 650 1160 670
<< locali >>
rect 965 1355 1215 1375
rect 965 1310 1215 1330
rect 965 765 1215 785
rect 90 670 115 765
rect 940 700 1105 720
rect 90 660 130 670
rect 90 640 100 660
rect 120 640 130 660
rect 90 630 130 640
rect 1085 610 1105 700
rect 1130 680 1150 765
rect 1130 670 1170 680
rect 1130 650 1140 670
rect 1160 650 1170 670
rect 1130 640 1170 650
<< metal1 >>
rect 990 1190 1215 1270
rect 990 1160 1045 1190
rect 1075 1160 1215 1190
rect 990 1080 1215 1160
rect 1010 935 1215 1015
rect 1010 905 1045 935
rect 1075 905 1215 935
rect 1010 825 1215 905
rect 715 695 795 710
rect 715 665 740 695
rect 770 665 795 695
rect 715 610 795 665
rect 1200 420 1215 610
rect 30 320 60 325
rect 30 295 40 320
rect 1200 165 1215 355
<< via1 >>
rect 1045 1160 1075 1190
rect 1045 905 1075 935
rect 740 665 770 695
rect 40 290 70 320
<< metal2 >>
rect 715 1190 1130 1265
rect 715 1160 1045 1190
rect 1075 1160 1130 1190
rect 715 1085 1130 1160
rect 715 695 795 1085
rect 715 665 740 695
rect 770 665 795 695
rect 715 645 795 665
rect 995 935 1130 1010
rect 995 905 1045 935
rect 1075 905 1130 935
rect 995 350 1130 905
rect 0 320 1130 350
rect 0 290 40 320
rect 70 290 1130 320
rect 0 265 1130 290
use dff_lower  dff_lower_0
timestamp 1620577227
transform 1 0 -35 0 1 130
box 30 -200 1250 505
use dff_upper  dff_upper_0
timestamp 1620577227
transform 1 0 -5 0 1 700
box 0 0 1015 695
<< labels >>
rlabel space -5 5 -5 5 7 clear
rlabel space -5 1365 -5 1365 7 preset
rlabel space -5 1320 -5 1320 7 CLK
rlabel space -5 775 -5 775 7 D
rlabel space -5 1175 -5 1175 7 VDD
rlabel space -5 920 -5 920 7 GND
rlabel locali 1215 775 1215 775 3 Q
<< end >>
