magic
tech sky130A
magscale 1 2
timestamp 1620712167
<< pwell >>
rect -4000 1643 -3204 1796
rect -4000 1153 -3847 1643
rect -3357 1153 -3204 1643
rect -4000 1000 -3204 1153
rect -3000 1643 -2204 1796
rect -3000 1153 -2847 1643
rect -2357 1153 -2204 1643
rect -3000 1000 -2204 1153
rect -2000 1643 -1204 1796
rect -2000 1153 -1847 1643
rect -1357 1153 -1204 1643
rect -2000 1000 -1204 1153
rect -1000 1643 -204 1796
rect -1000 1153 -847 1643
rect -357 1153 -204 1643
rect -1000 1000 -204 1153
rect 0 1643 796 1796
rect 0 1153 153 1643
rect 643 1153 796 1643
rect 0 1000 796 1153
rect 1000 1643 1796 1796
rect 1000 1153 1153 1643
rect 1643 1153 1796 1643
rect 1000 1000 1796 1153
rect -4000 643 -3204 796
rect -4000 153 -3847 643
rect -3357 153 -3204 643
rect -4000 0 -3204 153
rect -3000 643 -2204 796
rect -3000 153 -2847 643
rect -2357 153 -2204 643
rect -3000 0 -2204 153
rect -2000 643 -1204 796
rect -2000 153 -1847 643
rect -1357 153 -1204 643
rect -2000 0 -1204 153
rect -1000 643 -204 796
rect -1000 153 -847 643
rect -357 153 -204 643
rect -1000 0 -204 153
rect 0 643 796 796
rect 0 153 153 643
rect 643 153 796 643
rect 0 0 796 153
rect 1000 643 1796 796
rect 1000 153 1153 643
rect 1643 153 1796 643
rect 1000 0 1796 153
rect -4000 -357 -3204 -204
rect -4000 -847 -3847 -357
rect -3357 -847 -3204 -357
rect -4000 -1000 -3204 -847
rect -3000 -357 -2204 -204
rect -3000 -847 -2847 -357
rect -2357 -847 -2204 -357
rect -3000 -1000 -2204 -847
rect -2000 -357 -1204 -204
rect -2000 -847 -1847 -357
rect -1357 -847 -1204 -357
rect -2000 -1000 -1204 -847
rect -1000 -357 -204 -204
rect -1000 -847 -847 -357
rect -357 -847 -204 -357
rect -1000 -1000 -204 -847
rect 0 -357 796 -204
rect 0 -847 153 -357
rect 643 -847 796 -357
rect 0 -1000 796 -847
rect 1000 -357 1796 -204
rect 1000 -847 1153 -357
rect 1643 -847 1796 -357
rect 1000 -1000 1796 -847
rect -4000 -1357 -3204 -1204
rect -4000 -1847 -3847 -1357
rect -3357 -1847 -3204 -1357
rect -4000 -2000 -3204 -1847
rect -3000 -1357 -2204 -1204
rect -3000 -1847 -2847 -1357
rect -2357 -1847 -2204 -1357
rect -3000 -2000 -2204 -1847
rect -2000 -1357 -1204 -1204
rect -2000 -1847 -1847 -1357
rect -1357 -1847 -1204 -1357
rect -2000 -2000 -1204 -1847
rect -1000 -1357 -204 -1204
rect -1000 -1847 -847 -1357
rect -357 -1847 -204 -1357
rect -1000 -2000 -204 -1847
rect 0 -1357 796 -1204
rect 0 -1847 153 -1357
rect 643 -1847 796 -1357
rect 0 -2000 796 -1847
rect 1000 -1357 1796 -1204
rect 1000 -1847 1153 -1357
rect 1643 -1847 1796 -1357
rect 1000 -2000 1796 -1847
rect -4000 -2357 -3204 -2204
rect -4000 -2847 -3847 -2357
rect -3357 -2847 -3204 -2357
rect -4000 -3000 -3204 -2847
rect -3000 -2357 -2204 -2204
rect -3000 -2847 -2847 -2357
rect -2357 -2847 -2204 -2357
rect -3000 -3000 -2204 -2847
rect -2000 -2357 -1204 -2204
rect -2000 -2847 -1847 -2357
rect -1357 -2847 -1204 -2357
rect -2000 -3000 -1204 -2847
rect -1000 -2357 -204 -2204
rect -1000 -2847 -847 -2357
rect -357 -2847 -204 -2357
rect -1000 -3000 -204 -2847
rect 0 -2357 796 -2204
rect 0 -2847 153 -2357
rect 643 -2847 796 -2357
rect 0 -3000 796 -2847
rect 1000 -2357 1796 -2204
rect 1000 -2847 1153 -2357
rect 1643 -2847 1796 -2357
rect 1000 -3000 1796 -2847
<< nbase >>
rect -3847 1153 -3357 1643
rect -2847 1153 -2357 1643
rect -1847 1153 -1357 1643
rect -847 1153 -357 1643
rect 153 1153 643 1643
rect 1153 1153 1643 1643
rect -3847 153 -3357 643
rect -2847 153 -2357 643
rect -1847 153 -1357 643
rect -847 153 -357 643
rect 153 153 643 643
rect 1153 153 1643 643
rect -3847 -847 -3357 -357
rect -2847 -847 -2357 -357
rect -1847 -847 -1357 -357
rect -847 -847 -357 -357
rect 153 -847 643 -357
rect 1153 -847 1643 -357
rect -3847 -1847 -3357 -1357
rect -2847 -1847 -2357 -1357
rect -1847 -1847 -1357 -1357
rect -847 -1847 -357 -1357
rect 153 -1847 643 -1357
rect 1153 -1847 1643 -1357
rect -3847 -2847 -3357 -2357
rect -2847 -2847 -2357 -2357
rect -1847 -2847 -1357 -2357
rect -847 -2847 -357 -2357
rect 153 -2847 643 -2357
rect 1153 -2847 1643 -2357
<< pdiff >>
rect -3670 1449 -3534 1466
rect -3670 1347 -3653 1449
rect -3551 1347 -3534 1449
rect -3670 1330 -3534 1347
rect -2670 1449 -2534 1466
rect -2670 1347 -2653 1449
rect -2551 1347 -2534 1449
rect -2670 1330 -2534 1347
rect -1670 1449 -1534 1466
rect -1670 1347 -1653 1449
rect -1551 1347 -1534 1449
rect -1670 1330 -1534 1347
rect -670 1449 -534 1466
rect -670 1347 -653 1449
rect -551 1347 -534 1449
rect -670 1330 -534 1347
rect 330 1449 466 1466
rect 330 1347 347 1449
rect 449 1347 466 1449
rect 330 1330 466 1347
rect 1330 1449 1466 1466
rect 1330 1347 1347 1449
rect 1449 1347 1466 1449
rect 1330 1330 1466 1347
rect -3670 449 -3534 466
rect -3670 347 -3653 449
rect -3551 347 -3534 449
rect -3670 330 -3534 347
rect -2670 449 -2534 466
rect -2670 347 -2653 449
rect -2551 347 -2534 449
rect -2670 330 -2534 347
rect -1670 449 -1534 466
rect -1670 347 -1653 449
rect -1551 347 -1534 449
rect -1670 330 -1534 347
rect -670 449 -534 466
rect -670 347 -653 449
rect -551 347 -534 449
rect -670 330 -534 347
rect 330 449 466 466
rect 330 347 347 449
rect 449 347 466 449
rect 330 330 466 347
rect 1330 449 1466 466
rect 1330 347 1347 449
rect 1449 347 1466 449
rect 1330 330 1466 347
rect -3670 -551 -3534 -534
rect -3670 -653 -3653 -551
rect -3551 -653 -3534 -551
rect -3670 -670 -3534 -653
rect -2670 -551 -2534 -534
rect -2670 -653 -2653 -551
rect -2551 -653 -2534 -551
rect -2670 -670 -2534 -653
rect -1670 -551 -1534 -534
rect -1670 -653 -1653 -551
rect -1551 -653 -1534 -551
rect -1670 -670 -1534 -653
rect -670 -551 -534 -534
rect -670 -653 -653 -551
rect -551 -653 -534 -551
rect -670 -670 -534 -653
rect 330 -551 466 -534
rect 330 -653 347 -551
rect 449 -653 466 -551
rect 330 -670 466 -653
rect 1330 -551 1466 -534
rect 1330 -653 1347 -551
rect 1449 -653 1466 -551
rect 1330 -670 1466 -653
rect -3670 -1551 -3534 -1534
rect -3670 -1653 -3653 -1551
rect -3551 -1653 -3534 -1551
rect -3670 -1670 -3534 -1653
rect -2670 -1551 -2534 -1534
rect -2670 -1653 -2653 -1551
rect -2551 -1653 -2534 -1551
rect -2670 -1670 -2534 -1653
rect -1670 -1551 -1534 -1534
rect -1670 -1653 -1653 -1551
rect -1551 -1653 -1534 -1551
rect -1670 -1670 -1534 -1653
rect -670 -1551 -534 -1534
rect -670 -1653 -653 -1551
rect -551 -1653 -534 -1551
rect -670 -1670 -534 -1653
rect 330 -1551 466 -1534
rect 330 -1653 347 -1551
rect 449 -1653 466 -1551
rect 330 -1670 466 -1653
rect 1330 -1551 1466 -1534
rect 1330 -1653 1347 -1551
rect 1449 -1653 1466 -1551
rect 1330 -1670 1466 -1653
rect -3670 -2551 -3534 -2534
rect -3670 -2653 -3653 -2551
rect -3551 -2653 -3534 -2551
rect -3670 -2670 -3534 -2653
rect -2670 -2551 -2534 -2534
rect -2670 -2653 -2653 -2551
rect -2551 -2653 -2534 -2551
rect -2670 -2670 -2534 -2653
rect -1670 -2551 -1534 -2534
rect -1670 -2653 -1653 -2551
rect -1551 -2653 -1534 -2551
rect -1670 -2670 -1534 -2653
rect -670 -2551 -534 -2534
rect -670 -2653 -653 -2551
rect -551 -2653 -534 -2551
rect -670 -2670 -534 -2653
rect 330 -2551 466 -2534
rect 330 -2653 347 -2551
rect 449 -2653 466 -2551
rect 330 -2670 466 -2653
rect 1330 -2551 1466 -2534
rect 1330 -2653 1347 -2551
rect 1449 -2653 1466 -2551
rect 1330 -2670 1466 -2653
<< pdiffc >>
rect -3653 1347 -3551 1449
rect -2653 1347 -2551 1449
rect -1653 1347 -1551 1449
rect -653 1347 -551 1449
rect 347 1347 449 1449
rect 1347 1347 1449 1449
rect -3653 347 -3551 449
rect -2653 347 -2551 449
rect -1653 347 -1551 449
rect -653 347 -551 449
rect 347 347 449 449
rect 1347 347 1449 449
rect -3653 -653 -3551 -551
rect -2653 -653 -2551 -551
rect -1653 -653 -1551 -551
rect -653 -653 -551 -551
rect 347 -653 449 -551
rect 1347 -653 1449 -551
rect -3653 -1653 -3551 -1551
rect -2653 -1653 -2551 -1551
rect -1653 -1653 -1551 -1551
rect -653 -1653 -551 -1551
rect 347 -1653 449 -1551
rect 1347 -1653 1449 -1551
rect -3653 -2653 -3551 -2551
rect -2653 -2653 -2551 -2551
rect -1653 -2653 -1551 -2551
rect -653 -2653 -551 -2551
rect 347 -2653 449 -2551
rect 1347 -2653 1449 -2551
<< psubdiff >>
rect -3974 1736 -3230 1770
rect -3974 1702 -3940 1736
rect -3906 1702 -3872 1736
rect -3838 1702 -3804 1736
rect -3770 1702 -3736 1736
rect -3702 1702 -3502 1736
rect -3468 1702 -3434 1736
rect -3400 1702 -3366 1736
rect -3332 1702 -3298 1736
rect -3264 1702 -3230 1736
rect -3974 1669 -3230 1702
rect -3974 1668 -3873 1669
rect -3974 1634 -3940 1668
rect -3906 1634 -3873 1668
rect -3974 1600 -3873 1634
rect -3331 1668 -3230 1669
rect -3331 1634 -3298 1668
rect -3264 1634 -3230 1668
rect -3974 1566 -3940 1600
rect -3906 1566 -3873 1600
rect -3974 1532 -3873 1566
rect -3974 1498 -3940 1532
rect -3906 1498 -3873 1532
rect -3974 1298 -3873 1498
rect -3974 1264 -3940 1298
rect -3906 1264 -3873 1298
rect -3974 1230 -3873 1264
rect -3974 1196 -3940 1230
rect -3906 1196 -3873 1230
rect -3974 1162 -3873 1196
rect -3331 1600 -3230 1634
rect -3331 1566 -3298 1600
rect -3264 1566 -3230 1600
rect -3331 1532 -3230 1566
rect -3331 1498 -3298 1532
rect -3264 1498 -3230 1532
rect -3331 1298 -3230 1498
rect -3331 1264 -3298 1298
rect -3264 1264 -3230 1298
rect -3331 1230 -3230 1264
rect -3331 1196 -3298 1230
rect -3264 1196 -3230 1230
rect -3974 1128 -3940 1162
rect -3906 1128 -3873 1162
rect -3974 1127 -3873 1128
rect -3331 1162 -3230 1196
rect -3331 1128 -3298 1162
rect -3264 1128 -3230 1162
rect -3331 1127 -3230 1128
rect -3974 1094 -3230 1127
rect -3974 1060 -3940 1094
rect -3906 1060 -3872 1094
rect -3838 1060 -3804 1094
rect -3770 1060 -3736 1094
rect -3702 1060 -3502 1094
rect -3468 1060 -3434 1094
rect -3400 1060 -3366 1094
rect -3332 1060 -3298 1094
rect -3264 1060 -3230 1094
rect -3974 1026 -3230 1060
rect -2974 1736 -2230 1770
rect -2974 1702 -2940 1736
rect -2906 1702 -2872 1736
rect -2838 1702 -2804 1736
rect -2770 1702 -2736 1736
rect -2702 1702 -2502 1736
rect -2468 1702 -2434 1736
rect -2400 1702 -2366 1736
rect -2332 1702 -2298 1736
rect -2264 1702 -2230 1736
rect -2974 1669 -2230 1702
rect -2974 1668 -2873 1669
rect -2974 1634 -2940 1668
rect -2906 1634 -2873 1668
rect -2974 1600 -2873 1634
rect -2331 1668 -2230 1669
rect -2331 1634 -2298 1668
rect -2264 1634 -2230 1668
rect -2974 1566 -2940 1600
rect -2906 1566 -2873 1600
rect -2974 1532 -2873 1566
rect -2974 1498 -2940 1532
rect -2906 1498 -2873 1532
rect -2974 1298 -2873 1498
rect -2974 1264 -2940 1298
rect -2906 1264 -2873 1298
rect -2974 1230 -2873 1264
rect -2974 1196 -2940 1230
rect -2906 1196 -2873 1230
rect -2974 1162 -2873 1196
rect -2331 1600 -2230 1634
rect -2331 1566 -2298 1600
rect -2264 1566 -2230 1600
rect -2331 1532 -2230 1566
rect -2331 1498 -2298 1532
rect -2264 1498 -2230 1532
rect -2331 1298 -2230 1498
rect -2331 1264 -2298 1298
rect -2264 1264 -2230 1298
rect -2331 1230 -2230 1264
rect -2331 1196 -2298 1230
rect -2264 1196 -2230 1230
rect -2974 1128 -2940 1162
rect -2906 1128 -2873 1162
rect -2974 1127 -2873 1128
rect -2331 1162 -2230 1196
rect -2331 1128 -2298 1162
rect -2264 1128 -2230 1162
rect -2331 1127 -2230 1128
rect -2974 1094 -2230 1127
rect -2974 1060 -2940 1094
rect -2906 1060 -2872 1094
rect -2838 1060 -2804 1094
rect -2770 1060 -2736 1094
rect -2702 1060 -2502 1094
rect -2468 1060 -2434 1094
rect -2400 1060 -2366 1094
rect -2332 1060 -2298 1094
rect -2264 1060 -2230 1094
rect -2974 1026 -2230 1060
rect -1974 1736 -1230 1770
rect -1974 1702 -1940 1736
rect -1906 1702 -1872 1736
rect -1838 1702 -1804 1736
rect -1770 1702 -1736 1736
rect -1702 1702 -1502 1736
rect -1468 1702 -1434 1736
rect -1400 1702 -1366 1736
rect -1332 1702 -1298 1736
rect -1264 1702 -1230 1736
rect -1974 1669 -1230 1702
rect -1974 1668 -1873 1669
rect -1974 1634 -1940 1668
rect -1906 1634 -1873 1668
rect -1974 1600 -1873 1634
rect -1331 1668 -1230 1669
rect -1331 1634 -1298 1668
rect -1264 1634 -1230 1668
rect -1974 1566 -1940 1600
rect -1906 1566 -1873 1600
rect -1974 1532 -1873 1566
rect -1974 1498 -1940 1532
rect -1906 1498 -1873 1532
rect -1974 1298 -1873 1498
rect -1974 1264 -1940 1298
rect -1906 1264 -1873 1298
rect -1974 1230 -1873 1264
rect -1974 1196 -1940 1230
rect -1906 1196 -1873 1230
rect -1974 1162 -1873 1196
rect -1331 1600 -1230 1634
rect -1331 1566 -1298 1600
rect -1264 1566 -1230 1600
rect -1331 1532 -1230 1566
rect -1331 1498 -1298 1532
rect -1264 1498 -1230 1532
rect -1331 1298 -1230 1498
rect -1331 1264 -1298 1298
rect -1264 1264 -1230 1298
rect -1331 1230 -1230 1264
rect -1331 1196 -1298 1230
rect -1264 1196 -1230 1230
rect -1974 1128 -1940 1162
rect -1906 1128 -1873 1162
rect -1974 1127 -1873 1128
rect -1331 1162 -1230 1196
rect -1331 1128 -1298 1162
rect -1264 1128 -1230 1162
rect -1331 1127 -1230 1128
rect -1974 1094 -1230 1127
rect -1974 1060 -1940 1094
rect -1906 1060 -1872 1094
rect -1838 1060 -1804 1094
rect -1770 1060 -1736 1094
rect -1702 1060 -1502 1094
rect -1468 1060 -1434 1094
rect -1400 1060 -1366 1094
rect -1332 1060 -1298 1094
rect -1264 1060 -1230 1094
rect -1974 1026 -1230 1060
rect -974 1736 -230 1770
rect -974 1702 -940 1736
rect -906 1702 -872 1736
rect -838 1702 -804 1736
rect -770 1702 -736 1736
rect -702 1702 -502 1736
rect -468 1702 -434 1736
rect -400 1702 -366 1736
rect -332 1702 -298 1736
rect -264 1702 -230 1736
rect -974 1669 -230 1702
rect -974 1668 -873 1669
rect -974 1634 -940 1668
rect -906 1634 -873 1668
rect -974 1600 -873 1634
rect -331 1668 -230 1669
rect -331 1634 -298 1668
rect -264 1634 -230 1668
rect -974 1566 -940 1600
rect -906 1566 -873 1600
rect -974 1532 -873 1566
rect -974 1498 -940 1532
rect -906 1498 -873 1532
rect -974 1298 -873 1498
rect -974 1264 -940 1298
rect -906 1264 -873 1298
rect -974 1230 -873 1264
rect -974 1196 -940 1230
rect -906 1196 -873 1230
rect -974 1162 -873 1196
rect -331 1600 -230 1634
rect -331 1566 -298 1600
rect -264 1566 -230 1600
rect -331 1532 -230 1566
rect -331 1498 -298 1532
rect -264 1498 -230 1532
rect -331 1298 -230 1498
rect -331 1264 -298 1298
rect -264 1264 -230 1298
rect -331 1230 -230 1264
rect -331 1196 -298 1230
rect -264 1196 -230 1230
rect -974 1128 -940 1162
rect -906 1128 -873 1162
rect -974 1127 -873 1128
rect -331 1162 -230 1196
rect -331 1128 -298 1162
rect -264 1128 -230 1162
rect -331 1127 -230 1128
rect -974 1094 -230 1127
rect -974 1060 -940 1094
rect -906 1060 -872 1094
rect -838 1060 -804 1094
rect -770 1060 -736 1094
rect -702 1060 -502 1094
rect -468 1060 -434 1094
rect -400 1060 -366 1094
rect -332 1060 -298 1094
rect -264 1060 -230 1094
rect -974 1026 -230 1060
rect 26 1736 770 1770
rect 26 1702 60 1736
rect 94 1702 128 1736
rect 162 1702 196 1736
rect 230 1702 264 1736
rect 298 1702 498 1736
rect 532 1702 566 1736
rect 600 1702 634 1736
rect 668 1702 702 1736
rect 736 1702 770 1736
rect 26 1669 770 1702
rect 26 1668 127 1669
rect 26 1634 60 1668
rect 94 1634 127 1668
rect 26 1600 127 1634
rect 669 1668 770 1669
rect 669 1634 702 1668
rect 736 1634 770 1668
rect 26 1566 60 1600
rect 94 1566 127 1600
rect 26 1532 127 1566
rect 26 1498 60 1532
rect 94 1498 127 1532
rect 26 1298 127 1498
rect 26 1264 60 1298
rect 94 1264 127 1298
rect 26 1230 127 1264
rect 26 1196 60 1230
rect 94 1196 127 1230
rect 26 1162 127 1196
rect 669 1600 770 1634
rect 669 1566 702 1600
rect 736 1566 770 1600
rect 669 1532 770 1566
rect 669 1498 702 1532
rect 736 1498 770 1532
rect 669 1298 770 1498
rect 669 1264 702 1298
rect 736 1264 770 1298
rect 669 1230 770 1264
rect 669 1196 702 1230
rect 736 1196 770 1230
rect 26 1128 60 1162
rect 94 1128 127 1162
rect 26 1127 127 1128
rect 669 1162 770 1196
rect 669 1128 702 1162
rect 736 1128 770 1162
rect 669 1127 770 1128
rect 26 1094 770 1127
rect 26 1060 60 1094
rect 94 1060 128 1094
rect 162 1060 196 1094
rect 230 1060 264 1094
rect 298 1060 498 1094
rect 532 1060 566 1094
rect 600 1060 634 1094
rect 668 1060 702 1094
rect 736 1060 770 1094
rect 26 1026 770 1060
rect 1026 1736 1770 1770
rect 1026 1702 1060 1736
rect 1094 1702 1128 1736
rect 1162 1702 1196 1736
rect 1230 1702 1264 1736
rect 1298 1702 1498 1736
rect 1532 1702 1566 1736
rect 1600 1702 1634 1736
rect 1668 1702 1702 1736
rect 1736 1702 1770 1736
rect 1026 1669 1770 1702
rect 1026 1668 1127 1669
rect 1026 1634 1060 1668
rect 1094 1634 1127 1668
rect 1026 1600 1127 1634
rect 1669 1668 1770 1669
rect 1669 1634 1702 1668
rect 1736 1634 1770 1668
rect 1026 1566 1060 1600
rect 1094 1566 1127 1600
rect 1026 1532 1127 1566
rect 1026 1498 1060 1532
rect 1094 1498 1127 1532
rect 1026 1298 1127 1498
rect 1026 1264 1060 1298
rect 1094 1264 1127 1298
rect 1026 1230 1127 1264
rect 1026 1196 1060 1230
rect 1094 1196 1127 1230
rect 1026 1162 1127 1196
rect 1669 1600 1770 1634
rect 1669 1566 1702 1600
rect 1736 1566 1770 1600
rect 1669 1532 1770 1566
rect 1669 1498 1702 1532
rect 1736 1498 1770 1532
rect 1669 1298 1770 1498
rect 1669 1264 1702 1298
rect 1736 1264 1770 1298
rect 1669 1230 1770 1264
rect 1669 1196 1702 1230
rect 1736 1196 1770 1230
rect 1026 1128 1060 1162
rect 1094 1128 1127 1162
rect 1026 1127 1127 1128
rect 1669 1162 1770 1196
rect 1669 1128 1702 1162
rect 1736 1128 1770 1162
rect 1669 1127 1770 1128
rect 1026 1094 1770 1127
rect 1026 1060 1060 1094
rect 1094 1060 1128 1094
rect 1162 1060 1196 1094
rect 1230 1060 1264 1094
rect 1298 1060 1498 1094
rect 1532 1060 1566 1094
rect 1600 1060 1634 1094
rect 1668 1060 1702 1094
rect 1736 1060 1770 1094
rect 1026 1026 1770 1060
rect -3974 736 -3230 770
rect -3974 702 -3940 736
rect -3906 702 -3872 736
rect -3838 702 -3804 736
rect -3770 702 -3736 736
rect -3702 702 -3502 736
rect -3468 702 -3434 736
rect -3400 702 -3366 736
rect -3332 702 -3298 736
rect -3264 702 -3230 736
rect -3974 669 -3230 702
rect -3974 668 -3873 669
rect -3974 634 -3940 668
rect -3906 634 -3873 668
rect -3974 600 -3873 634
rect -3331 668 -3230 669
rect -3331 634 -3298 668
rect -3264 634 -3230 668
rect -3974 566 -3940 600
rect -3906 566 -3873 600
rect -3974 532 -3873 566
rect -3974 498 -3940 532
rect -3906 498 -3873 532
rect -3974 298 -3873 498
rect -3974 264 -3940 298
rect -3906 264 -3873 298
rect -3974 230 -3873 264
rect -3974 196 -3940 230
rect -3906 196 -3873 230
rect -3974 162 -3873 196
rect -3331 600 -3230 634
rect -3331 566 -3298 600
rect -3264 566 -3230 600
rect -3331 532 -3230 566
rect -3331 498 -3298 532
rect -3264 498 -3230 532
rect -3331 298 -3230 498
rect -3331 264 -3298 298
rect -3264 264 -3230 298
rect -3331 230 -3230 264
rect -3331 196 -3298 230
rect -3264 196 -3230 230
rect -3974 128 -3940 162
rect -3906 128 -3873 162
rect -3974 127 -3873 128
rect -3331 162 -3230 196
rect -3331 128 -3298 162
rect -3264 128 -3230 162
rect -3331 127 -3230 128
rect -3974 94 -3230 127
rect -3974 60 -3940 94
rect -3906 60 -3872 94
rect -3838 60 -3804 94
rect -3770 60 -3736 94
rect -3702 60 -3502 94
rect -3468 60 -3434 94
rect -3400 60 -3366 94
rect -3332 60 -3298 94
rect -3264 60 -3230 94
rect -3974 26 -3230 60
rect -2974 736 -2230 770
rect -2974 702 -2940 736
rect -2906 702 -2872 736
rect -2838 702 -2804 736
rect -2770 702 -2736 736
rect -2702 702 -2502 736
rect -2468 702 -2434 736
rect -2400 702 -2366 736
rect -2332 702 -2298 736
rect -2264 702 -2230 736
rect -2974 669 -2230 702
rect -2974 668 -2873 669
rect -2974 634 -2940 668
rect -2906 634 -2873 668
rect -2974 600 -2873 634
rect -2331 668 -2230 669
rect -2331 634 -2298 668
rect -2264 634 -2230 668
rect -2974 566 -2940 600
rect -2906 566 -2873 600
rect -2974 532 -2873 566
rect -2974 498 -2940 532
rect -2906 498 -2873 532
rect -2974 298 -2873 498
rect -2974 264 -2940 298
rect -2906 264 -2873 298
rect -2974 230 -2873 264
rect -2974 196 -2940 230
rect -2906 196 -2873 230
rect -2974 162 -2873 196
rect -2331 600 -2230 634
rect -2331 566 -2298 600
rect -2264 566 -2230 600
rect -2331 532 -2230 566
rect -2331 498 -2298 532
rect -2264 498 -2230 532
rect -2331 298 -2230 498
rect -2331 264 -2298 298
rect -2264 264 -2230 298
rect -2331 230 -2230 264
rect -2331 196 -2298 230
rect -2264 196 -2230 230
rect -2974 128 -2940 162
rect -2906 128 -2873 162
rect -2974 127 -2873 128
rect -2331 162 -2230 196
rect -2331 128 -2298 162
rect -2264 128 -2230 162
rect -2331 127 -2230 128
rect -2974 94 -2230 127
rect -2974 60 -2940 94
rect -2906 60 -2872 94
rect -2838 60 -2804 94
rect -2770 60 -2736 94
rect -2702 60 -2502 94
rect -2468 60 -2434 94
rect -2400 60 -2366 94
rect -2332 60 -2298 94
rect -2264 60 -2230 94
rect -2974 26 -2230 60
rect -1974 736 -1230 770
rect -1974 702 -1940 736
rect -1906 702 -1872 736
rect -1838 702 -1804 736
rect -1770 702 -1736 736
rect -1702 702 -1502 736
rect -1468 702 -1434 736
rect -1400 702 -1366 736
rect -1332 702 -1298 736
rect -1264 702 -1230 736
rect -1974 669 -1230 702
rect -1974 668 -1873 669
rect -1974 634 -1940 668
rect -1906 634 -1873 668
rect -1974 600 -1873 634
rect -1331 668 -1230 669
rect -1331 634 -1298 668
rect -1264 634 -1230 668
rect -1974 566 -1940 600
rect -1906 566 -1873 600
rect -1974 532 -1873 566
rect -1974 498 -1940 532
rect -1906 498 -1873 532
rect -1974 298 -1873 498
rect -1974 264 -1940 298
rect -1906 264 -1873 298
rect -1974 230 -1873 264
rect -1974 196 -1940 230
rect -1906 196 -1873 230
rect -1974 162 -1873 196
rect -1331 600 -1230 634
rect -1331 566 -1298 600
rect -1264 566 -1230 600
rect -1331 532 -1230 566
rect -1331 498 -1298 532
rect -1264 498 -1230 532
rect -1331 298 -1230 498
rect -1331 264 -1298 298
rect -1264 264 -1230 298
rect -1331 230 -1230 264
rect -1331 196 -1298 230
rect -1264 196 -1230 230
rect -1974 128 -1940 162
rect -1906 128 -1873 162
rect -1974 127 -1873 128
rect -1331 162 -1230 196
rect -1331 128 -1298 162
rect -1264 128 -1230 162
rect -1331 127 -1230 128
rect -1974 94 -1230 127
rect -1974 60 -1940 94
rect -1906 60 -1872 94
rect -1838 60 -1804 94
rect -1770 60 -1736 94
rect -1702 60 -1502 94
rect -1468 60 -1434 94
rect -1400 60 -1366 94
rect -1332 60 -1298 94
rect -1264 60 -1230 94
rect -1974 26 -1230 60
rect -974 736 -230 770
rect -974 702 -940 736
rect -906 702 -872 736
rect -838 702 -804 736
rect -770 702 -736 736
rect -702 702 -502 736
rect -468 702 -434 736
rect -400 702 -366 736
rect -332 702 -298 736
rect -264 702 -230 736
rect -974 669 -230 702
rect -974 668 -873 669
rect -974 634 -940 668
rect -906 634 -873 668
rect -974 600 -873 634
rect -331 668 -230 669
rect -331 634 -298 668
rect -264 634 -230 668
rect -974 566 -940 600
rect -906 566 -873 600
rect -974 532 -873 566
rect -974 498 -940 532
rect -906 498 -873 532
rect -974 298 -873 498
rect -974 264 -940 298
rect -906 264 -873 298
rect -974 230 -873 264
rect -974 196 -940 230
rect -906 196 -873 230
rect -974 162 -873 196
rect -331 600 -230 634
rect -331 566 -298 600
rect -264 566 -230 600
rect -331 532 -230 566
rect -331 498 -298 532
rect -264 498 -230 532
rect -331 298 -230 498
rect -331 264 -298 298
rect -264 264 -230 298
rect -331 230 -230 264
rect -331 196 -298 230
rect -264 196 -230 230
rect -974 128 -940 162
rect -906 128 -873 162
rect -974 127 -873 128
rect -331 162 -230 196
rect -331 128 -298 162
rect -264 128 -230 162
rect -331 127 -230 128
rect -974 94 -230 127
rect -974 60 -940 94
rect -906 60 -872 94
rect -838 60 -804 94
rect -770 60 -736 94
rect -702 60 -502 94
rect -468 60 -434 94
rect -400 60 -366 94
rect -332 60 -298 94
rect -264 60 -230 94
rect -974 26 -230 60
rect 26 736 770 770
rect 26 702 60 736
rect 94 702 128 736
rect 162 702 196 736
rect 230 702 264 736
rect 298 702 498 736
rect 532 702 566 736
rect 600 702 634 736
rect 668 702 702 736
rect 736 702 770 736
rect 26 669 770 702
rect 26 668 127 669
rect 26 634 60 668
rect 94 634 127 668
rect 26 600 127 634
rect 669 668 770 669
rect 669 634 702 668
rect 736 634 770 668
rect 26 566 60 600
rect 94 566 127 600
rect 26 532 127 566
rect 26 498 60 532
rect 94 498 127 532
rect 26 298 127 498
rect 26 264 60 298
rect 94 264 127 298
rect 26 230 127 264
rect 26 196 60 230
rect 94 196 127 230
rect 26 162 127 196
rect 669 600 770 634
rect 669 566 702 600
rect 736 566 770 600
rect 669 532 770 566
rect 669 498 702 532
rect 736 498 770 532
rect 669 298 770 498
rect 669 264 702 298
rect 736 264 770 298
rect 669 230 770 264
rect 669 196 702 230
rect 736 196 770 230
rect 26 128 60 162
rect 94 128 127 162
rect 26 127 127 128
rect 669 162 770 196
rect 669 128 702 162
rect 736 128 770 162
rect 669 127 770 128
rect 26 94 770 127
rect 26 60 60 94
rect 94 60 128 94
rect 162 60 196 94
rect 230 60 264 94
rect 298 60 498 94
rect 532 60 566 94
rect 600 60 634 94
rect 668 60 702 94
rect 736 60 770 94
rect 26 26 770 60
rect 1026 736 1770 770
rect 1026 702 1060 736
rect 1094 702 1128 736
rect 1162 702 1196 736
rect 1230 702 1264 736
rect 1298 702 1498 736
rect 1532 702 1566 736
rect 1600 702 1634 736
rect 1668 702 1702 736
rect 1736 702 1770 736
rect 1026 669 1770 702
rect 1026 668 1127 669
rect 1026 634 1060 668
rect 1094 634 1127 668
rect 1026 600 1127 634
rect 1669 668 1770 669
rect 1669 634 1702 668
rect 1736 634 1770 668
rect 1026 566 1060 600
rect 1094 566 1127 600
rect 1026 532 1127 566
rect 1026 498 1060 532
rect 1094 498 1127 532
rect 1026 298 1127 498
rect 1026 264 1060 298
rect 1094 264 1127 298
rect 1026 230 1127 264
rect 1026 196 1060 230
rect 1094 196 1127 230
rect 1026 162 1127 196
rect 1669 600 1770 634
rect 1669 566 1702 600
rect 1736 566 1770 600
rect 1669 532 1770 566
rect 1669 498 1702 532
rect 1736 498 1770 532
rect 1669 298 1770 498
rect 1669 264 1702 298
rect 1736 264 1770 298
rect 1669 230 1770 264
rect 1669 196 1702 230
rect 1736 196 1770 230
rect 1026 128 1060 162
rect 1094 128 1127 162
rect 1026 127 1127 128
rect 1669 162 1770 196
rect 1669 128 1702 162
rect 1736 128 1770 162
rect 1669 127 1770 128
rect 1026 94 1770 127
rect 1026 60 1060 94
rect 1094 60 1128 94
rect 1162 60 1196 94
rect 1230 60 1264 94
rect 1298 60 1498 94
rect 1532 60 1566 94
rect 1600 60 1634 94
rect 1668 60 1702 94
rect 1736 60 1770 94
rect 1026 26 1770 60
rect -3974 -264 -3230 -230
rect -3974 -298 -3940 -264
rect -3906 -298 -3872 -264
rect -3838 -298 -3804 -264
rect -3770 -298 -3736 -264
rect -3702 -298 -3502 -264
rect -3468 -298 -3434 -264
rect -3400 -298 -3366 -264
rect -3332 -298 -3298 -264
rect -3264 -298 -3230 -264
rect -3974 -331 -3230 -298
rect -3974 -332 -3873 -331
rect -3974 -366 -3940 -332
rect -3906 -366 -3873 -332
rect -3974 -400 -3873 -366
rect -3331 -332 -3230 -331
rect -3331 -366 -3298 -332
rect -3264 -366 -3230 -332
rect -3974 -434 -3940 -400
rect -3906 -434 -3873 -400
rect -3974 -468 -3873 -434
rect -3974 -502 -3940 -468
rect -3906 -502 -3873 -468
rect -3974 -702 -3873 -502
rect -3974 -736 -3940 -702
rect -3906 -736 -3873 -702
rect -3974 -770 -3873 -736
rect -3974 -804 -3940 -770
rect -3906 -804 -3873 -770
rect -3974 -838 -3873 -804
rect -3331 -400 -3230 -366
rect -3331 -434 -3298 -400
rect -3264 -434 -3230 -400
rect -3331 -468 -3230 -434
rect -3331 -502 -3298 -468
rect -3264 -502 -3230 -468
rect -3331 -702 -3230 -502
rect -3331 -736 -3298 -702
rect -3264 -736 -3230 -702
rect -3331 -770 -3230 -736
rect -3331 -804 -3298 -770
rect -3264 -804 -3230 -770
rect -3974 -872 -3940 -838
rect -3906 -872 -3873 -838
rect -3974 -873 -3873 -872
rect -3331 -838 -3230 -804
rect -3331 -872 -3298 -838
rect -3264 -872 -3230 -838
rect -3331 -873 -3230 -872
rect -3974 -906 -3230 -873
rect -3974 -940 -3940 -906
rect -3906 -940 -3872 -906
rect -3838 -940 -3804 -906
rect -3770 -940 -3736 -906
rect -3702 -940 -3502 -906
rect -3468 -940 -3434 -906
rect -3400 -940 -3366 -906
rect -3332 -940 -3298 -906
rect -3264 -940 -3230 -906
rect -3974 -974 -3230 -940
rect -2974 -264 -2230 -230
rect -2974 -298 -2940 -264
rect -2906 -298 -2872 -264
rect -2838 -298 -2804 -264
rect -2770 -298 -2736 -264
rect -2702 -298 -2502 -264
rect -2468 -298 -2434 -264
rect -2400 -298 -2366 -264
rect -2332 -298 -2298 -264
rect -2264 -298 -2230 -264
rect -2974 -331 -2230 -298
rect -2974 -332 -2873 -331
rect -2974 -366 -2940 -332
rect -2906 -366 -2873 -332
rect -2974 -400 -2873 -366
rect -2331 -332 -2230 -331
rect -2331 -366 -2298 -332
rect -2264 -366 -2230 -332
rect -2974 -434 -2940 -400
rect -2906 -434 -2873 -400
rect -2974 -468 -2873 -434
rect -2974 -502 -2940 -468
rect -2906 -502 -2873 -468
rect -2974 -702 -2873 -502
rect -2974 -736 -2940 -702
rect -2906 -736 -2873 -702
rect -2974 -770 -2873 -736
rect -2974 -804 -2940 -770
rect -2906 -804 -2873 -770
rect -2974 -838 -2873 -804
rect -2331 -400 -2230 -366
rect -2331 -434 -2298 -400
rect -2264 -434 -2230 -400
rect -2331 -468 -2230 -434
rect -2331 -502 -2298 -468
rect -2264 -502 -2230 -468
rect -2331 -702 -2230 -502
rect -2331 -736 -2298 -702
rect -2264 -736 -2230 -702
rect -2331 -770 -2230 -736
rect -2331 -804 -2298 -770
rect -2264 -804 -2230 -770
rect -2974 -872 -2940 -838
rect -2906 -872 -2873 -838
rect -2974 -873 -2873 -872
rect -2331 -838 -2230 -804
rect -2331 -872 -2298 -838
rect -2264 -872 -2230 -838
rect -2331 -873 -2230 -872
rect -2974 -906 -2230 -873
rect -2974 -940 -2940 -906
rect -2906 -940 -2872 -906
rect -2838 -940 -2804 -906
rect -2770 -940 -2736 -906
rect -2702 -940 -2502 -906
rect -2468 -940 -2434 -906
rect -2400 -940 -2366 -906
rect -2332 -940 -2298 -906
rect -2264 -940 -2230 -906
rect -2974 -974 -2230 -940
rect -1974 -264 -1230 -230
rect -1974 -298 -1940 -264
rect -1906 -298 -1872 -264
rect -1838 -298 -1804 -264
rect -1770 -298 -1736 -264
rect -1702 -298 -1502 -264
rect -1468 -298 -1434 -264
rect -1400 -298 -1366 -264
rect -1332 -298 -1298 -264
rect -1264 -298 -1230 -264
rect -1974 -331 -1230 -298
rect -1974 -332 -1873 -331
rect -1974 -366 -1940 -332
rect -1906 -366 -1873 -332
rect -1974 -400 -1873 -366
rect -1331 -332 -1230 -331
rect -1331 -366 -1298 -332
rect -1264 -366 -1230 -332
rect -1974 -434 -1940 -400
rect -1906 -434 -1873 -400
rect -1974 -468 -1873 -434
rect -1974 -502 -1940 -468
rect -1906 -502 -1873 -468
rect -1974 -702 -1873 -502
rect -1974 -736 -1940 -702
rect -1906 -736 -1873 -702
rect -1974 -770 -1873 -736
rect -1974 -804 -1940 -770
rect -1906 -804 -1873 -770
rect -1974 -838 -1873 -804
rect -1331 -400 -1230 -366
rect -1331 -434 -1298 -400
rect -1264 -434 -1230 -400
rect -1331 -468 -1230 -434
rect -1331 -502 -1298 -468
rect -1264 -502 -1230 -468
rect -1331 -702 -1230 -502
rect -1331 -736 -1298 -702
rect -1264 -736 -1230 -702
rect -1331 -770 -1230 -736
rect -1331 -804 -1298 -770
rect -1264 -804 -1230 -770
rect -1974 -872 -1940 -838
rect -1906 -872 -1873 -838
rect -1974 -873 -1873 -872
rect -1331 -838 -1230 -804
rect -1331 -872 -1298 -838
rect -1264 -872 -1230 -838
rect -1331 -873 -1230 -872
rect -1974 -906 -1230 -873
rect -1974 -940 -1940 -906
rect -1906 -940 -1872 -906
rect -1838 -940 -1804 -906
rect -1770 -940 -1736 -906
rect -1702 -940 -1502 -906
rect -1468 -940 -1434 -906
rect -1400 -940 -1366 -906
rect -1332 -940 -1298 -906
rect -1264 -940 -1230 -906
rect -1974 -974 -1230 -940
rect -974 -264 -230 -230
rect -974 -298 -940 -264
rect -906 -298 -872 -264
rect -838 -298 -804 -264
rect -770 -298 -736 -264
rect -702 -298 -502 -264
rect -468 -298 -434 -264
rect -400 -298 -366 -264
rect -332 -298 -298 -264
rect -264 -298 -230 -264
rect -974 -331 -230 -298
rect -974 -332 -873 -331
rect -974 -366 -940 -332
rect -906 -366 -873 -332
rect -974 -400 -873 -366
rect -331 -332 -230 -331
rect -331 -366 -298 -332
rect -264 -366 -230 -332
rect -974 -434 -940 -400
rect -906 -434 -873 -400
rect -974 -468 -873 -434
rect -974 -502 -940 -468
rect -906 -502 -873 -468
rect -974 -702 -873 -502
rect -974 -736 -940 -702
rect -906 -736 -873 -702
rect -974 -770 -873 -736
rect -974 -804 -940 -770
rect -906 -804 -873 -770
rect -974 -838 -873 -804
rect -331 -400 -230 -366
rect -331 -434 -298 -400
rect -264 -434 -230 -400
rect -331 -468 -230 -434
rect -331 -502 -298 -468
rect -264 -502 -230 -468
rect -331 -702 -230 -502
rect -331 -736 -298 -702
rect -264 -736 -230 -702
rect -331 -770 -230 -736
rect -331 -804 -298 -770
rect -264 -804 -230 -770
rect -974 -872 -940 -838
rect -906 -872 -873 -838
rect -974 -873 -873 -872
rect -331 -838 -230 -804
rect -331 -872 -298 -838
rect -264 -872 -230 -838
rect -331 -873 -230 -872
rect -974 -906 -230 -873
rect -974 -940 -940 -906
rect -906 -940 -872 -906
rect -838 -940 -804 -906
rect -770 -940 -736 -906
rect -702 -940 -502 -906
rect -468 -940 -434 -906
rect -400 -940 -366 -906
rect -332 -940 -298 -906
rect -264 -940 -230 -906
rect -974 -974 -230 -940
rect 26 -264 770 -230
rect 26 -298 60 -264
rect 94 -298 128 -264
rect 162 -298 196 -264
rect 230 -298 264 -264
rect 298 -298 498 -264
rect 532 -298 566 -264
rect 600 -298 634 -264
rect 668 -298 702 -264
rect 736 -298 770 -264
rect 26 -331 770 -298
rect 26 -332 127 -331
rect 26 -366 60 -332
rect 94 -366 127 -332
rect 26 -400 127 -366
rect 669 -332 770 -331
rect 669 -366 702 -332
rect 736 -366 770 -332
rect 26 -434 60 -400
rect 94 -434 127 -400
rect 26 -468 127 -434
rect 26 -502 60 -468
rect 94 -502 127 -468
rect 26 -702 127 -502
rect 26 -736 60 -702
rect 94 -736 127 -702
rect 26 -770 127 -736
rect 26 -804 60 -770
rect 94 -804 127 -770
rect 26 -838 127 -804
rect 669 -400 770 -366
rect 669 -434 702 -400
rect 736 -434 770 -400
rect 669 -468 770 -434
rect 669 -502 702 -468
rect 736 -502 770 -468
rect 669 -702 770 -502
rect 669 -736 702 -702
rect 736 -736 770 -702
rect 669 -770 770 -736
rect 669 -804 702 -770
rect 736 -804 770 -770
rect 26 -872 60 -838
rect 94 -872 127 -838
rect 26 -873 127 -872
rect 669 -838 770 -804
rect 669 -872 702 -838
rect 736 -872 770 -838
rect 669 -873 770 -872
rect 26 -906 770 -873
rect 26 -940 60 -906
rect 94 -940 128 -906
rect 162 -940 196 -906
rect 230 -940 264 -906
rect 298 -940 498 -906
rect 532 -940 566 -906
rect 600 -940 634 -906
rect 668 -940 702 -906
rect 736 -940 770 -906
rect 26 -974 770 -940
rect 1026 -264 1770 -230
rect 1026 -298 1060 -264
rect 1094 -298 1128 -264
rect 1162 -298 1196 -264
rect 1230 -298 1264 -264
rect 1298 -298 1498 -264
rect 1532 -298 1566 -264
rect 1600 -298 1634 -264
rect 1668 -298 1702 -264
rect 1736 -298 1770 -264
rect 1026 -331 1770 -298
rect 1026 -332 1127 -331
rect 1026 -366 1060 -332
rect 1094 -366 1127 -332
rect 1026 -400 1127 -366
rect 1669 -332 1770 -331
rect 1669 -366 1702 -332
rect 1736 -366 1770 -332
rect 1026 -434 1060 -400
rect 1094 -434 1127 -400
rect 1026 -468 1127 -434
rect 1026 -502 1060 -468
rect 1094 -502 1127 -468
rect 1026 -702 1127 -502
rect 1026 -736 1060 -702
rect 1094 -736 1127 -702
rect 1026 -770 1127 -736
rect 1026 -804 1060 -770
rect 1094 -804 1127 -770
rect 1026 -838 1127 -804
rect 1669 -400 1770 -366
rect 1669 -434 1702 -400
rect 1736 -434 1770 -400
rect 1669 -468 1770 -434
rect 1669 -502 1702 -468
rect 1736 -502 1770 -468
rect 1669 -702 1770 -502
rect 1669 -736 1702 -702
rect 1736 -736 1770 -702
rect 1669 -770 1770 -736
rect 1669 -804 1702 -770
rect 1736 -804 1770 -770
rect 1026 -872 1060 -838
rect 1094 -872 1127 -838
rect 1026 -873 1127 -872
rect 1669 -838 1770 -804
rect 1669 -872 1702 -838
rect 1736 -872 1770 -838
rect 1669 -873 1770 -872
rect 1026 -906 1770 -873
rect 1026 -940 1060 -906
rect 1094 -940 1128 -906
rect 1162 -940 1196 -906
rect 1230 -940 1264 -906
rect 1298 -940 1498 -906
rect 1532 -940 1566 -906
rect 1600 -940 1634 -906
rect 1668 -940 1702 -906
rect 1736 -940 1770 -906
rect 1026 -974 1770 -940
rect -3974 -1264 -3230 -1230
rect -3974 -1298 -3940 -1264
rect -3906 -1298 -3872 -1264
rect -3838 -1298 -3804 -1264
rect -3770 -1298 -3736 -1264
rect -3702 -1298 -3502 -1264
rect -3468 -1298 -3434 -1264
rect -3400 -1298 -3366 -1264
rect -3332 -1298 -3298 -1264
rect -3264 -1298 -3230 -1264
rect -3974 -1331 -3230 -1298
rect -3974 -1332 -3873 -1331
rect -3974 -1366 -3940 -1332
rect -3906 -1366 -3873 -1332
rect -3974 -1400 -3873 -1366
rect -3331 -1332 -3230 -1331
rect -3331 -1366 -3298 -1332
rect -3264 -1366 -3230 -1332
rect -3974 -1434 -3940 -1400
rect -3906 -1434 -3873 -1400
rect -3974 -1468 -3873 -1434
rect -3974 -1502 -3940 -1468
rect -3906 -1502 -3873 -1468
rect -3974 -1702 -3873 -1502
rect -3974 -1736 -3940 -1702
rect -3906 -1736 -3873 -1702
rect -3974 -1770 -3873 -1736
rect -3974 -1804 -3940 -1770
rect -3906 -1804 -3873 -1770
rect -3974 -1838 -3873 -1804
rect -3331 -1400 -3230 -1366
rect -3331 -1434 -3298 -1400
rect -3264 -1434 -3230 -1400
rect -3331 -1468 -3230 -1434
rect -3331 -1502 -3298 -1468
rect -3264 -1502 -3230 -1468
rect -3331 -1702 -3230 -1502
rect -3331 -1736 -3298 -1702
rect -3264 -1736 -3230 -1702
rect -3331 -1770 -3230 -1736
rect -3331 -1804 -3298 -1770
rect -3264 -1804 -3230 -1770
rect -3974 -1872 -3940 -1838
rect -3906 -1872 -3873 -1838
rect -3974 -1873 -3873 -1872
rect -3331 -1838 -3230 -1804
rect -3331 -1872 -3298 -1838
rect -3264 -1872 -3230 -1838
rect -3331 -1873 -3230 -1872
rect -3974 -1906 -3230 -1873
rect -3974 -1940 -3940 -1906
rect -3906 -1940 -3872 -1906
rect -3838 -1940 -3804 -1906
rect -3770 -1940 -3736 -1906
rect -3702 -1940 -3502 -1906
rect -3468 -1940 -3434 -1906
rect -3400 -1940 -3366 -1906
rect -3332 -1940 -3298 -1906
rect -3264 -1940 -3230 -1906
rect -3974 -1974 -3230 -1940
rect -2974 -1264 -2230 -1230
rect -2974 -1298 -2940 -1264
rect -2906 -1298 -2872 -1264
rect -2838 -1298 -2804 -1264
rect -2770 -1298 -2736 -1264
rect -2702 -1298 -2502 -1264
rect -2468 -1298 -2434 -1264
rect -2400 -1298 -2366 -1264
rect -2332 -1298 -2298 -1264
rect -2264 -1298 -2230 -1264
rect -2974 -1331 -2230 -1298
rect -2974 -1332 -2873 -1331
rect -2974 -1366 -2940 -1332
rect -2906 -1366 -2873 -1332
rect -2974 -1400 -2873 -1366
rect -2331 -1332 -2230 -1331
rect -2331 -1366 -2298 -1332
rect -2264 -1366 -2230 -1332
rect -2974 -1434 -2940 -1400
rect -2906 -1434 -2873 -1400
rect -2974 -1468 -2873 -1434
rect -2974 -1502 -2940 -1468
rect -2906 -1502 -2873 -1468
rect -2974 -1702 -2873 -1502
rect -2974 -1736 -2940 -1702
rect -2906 -1736 -2873 -1702
rect -2974 -1770 -2873 -1736
rect -2974 -1804 -2940 -1770
rect -2906 -1804 -2873 -1770
rect -2974 -1838 -2873 -1804
rect -2331 -1400 -2230 -1366
rect -2331 -1434 -2298 -1400
rect -2264 -1434 -2230 -1400
rect -2331 -1468 -2230 -1434
rect -2331 -1502 -2298 -1468
rect -2264 -1502 -2230 -1468
rect -2331 -1702 -2230 -1502
rect -2331 -1736 -2298 -1702
rect -2264 -1736 -2230 -1702
rect -2331 -1770 -2230 -1736
rect -2331 -1804 -2298 -1770
rect -2264 -1804 -2230 -1770
rect -2974 -1872 -2940 -1838
rect -2906 -1872 -2873 -1838
rect -2974 -1873 -2873 -1872
rect -2331 -1838 -2230 -1804
rect -2331 -1872 -2298 -1838
rect -2264 -1872 -2230 -1838
rect -2331 -1873 -2230 -1872
rect -2974 -1906 -2230 -1873
rect -2974 -1940 -2940 -1906
rect -2906 -1940 -2872 -1906
rect -2838 -1940 -2804 -1906
rect -2770 -1940 -2736 -1906
rect -2702 -1940 -2502 -1906
rect -2468 -1940 -2434 -1906
rect -2400 -1940 -2366 -1906
rect -2332 -1940 -2298 -1906
rect -2264 -1940 -2230 -1906
rect -2974 -1974 -2230 -1940
rect -1974 -1264 -1230 -1230
rect -1974 -1298 -1940 -1264
rect -1906 -1298 -1872 -1264
rect -1838 -1298 -1804 -1264
rect -1770 -1298 -1736 -1264
rect -1702 -1298 -1502 -1264
rect -1468 -1298 -1434 -1264
rect -1400 -1298 -1366 -1264
rect -1332 -1298 -1298 -1264
rect -1264 -1298 -1230 -1264
rect -1974 -1331 -1230 -1298
rect -1974 -1332 -1873 -1331
rect -1974 -1366 -1940 -1332
rect -1906 -1366 -1873 -1332
rect -1974 -1400 -1873 -1366
rect -1331 -1332 -1230 -1331
rect -1331 -1366 -1298 -1332
rect -1264 -1366 -1230 -1332
rect -1974 -1434 -1940 -1400
rect -1906 -1434 -1873 -1400
rect -1974 -1468 -1873 -1434
rect -1974 -1502 -1940 -1468
rect -1906 -1502 -1873 -1468
rect -1974 -1702 -1873 -1502
rect -1974 -1736 -1940 -1702
rect -1906 -1736 -1873 -1702
rect -1974 -1770 -1873 -1736
rect -1974 -1804 -1940 -1770
rect -1906 -1804 -1873 -1770
rect -1974 -1838 -1873 -1804
rect -1331 -1400 -1230 -1366
rect -1331 -1434 -1298 -1400
rect -1264 -1434 -1230 -1400
rect -1331 -1468 -1230 -1434
rect -1331 -1502 -1298 -1468
rect -1264 -1502 -1230 -1468
rect -1331 -1702 -1230 -1502
rect -1331 -1736 -1298 -1702
rect -1264 -1736 -1230 -1702
rect -1331 -1770 -1230 -1736
rect -1331 -1804 -1298 -1770
rect -1264 -1804 -1230 -1770
rect -1974 -1872 -1940 -1838
rect -1906 -1872 -1873 -1838
rect -1974 -1873 -1873 -1872
rect -1331 -1838 -1230 -1804
rect -1331 -1872 -1298 -1838
rect -1264 -1872 -1230 -1838
rect -1331 -1873 -1230 -1872
rect -1974 -1906 -1230 -1873
rect -1974 -1940 -1940 -1906
rect -1906 -1940 -1872 -1906
rect -1838 -1940 -1804 -1906
rect -1770 -1940 -1736 -1906
rect -1702 -1940 -1502 -1906
rect -1468 -1940 -1434 -1906
rect -1400 -1940 -1366 -1906
rect -1332 -1940 -1298 -1906
rect -1264 -1940 -1230 -1906
rect -1974 -1974 -1230 -1940
rect -974 -1264 -230 -1230
rect -974 -1298 -940 -1264
rect -906 -1298 -872 -1264
rect -838 -1298 -804 -1264
rect -770 -1298 -736 -1264
rect -702 -1298 -502 -1264
rect -468 -1298 -434 -1264
rect -400 -1298 -366 -1264
rect -332 -1298 -298 -1264
rect -264 -1298 -230 -1264
rect -974 -1331 -230 -1298
rect -974 -1332 -873 -1331
rect -974 -1366 -940 -1332
rect -906 -1366 -873 -1332
rect -974 -1400 -873 -1366
rect -331 -1332 -230 -1331
rect -331 -1366 -298 -1332
rect -264 -1366 -230 -1332
rect -974 -1434 -940 -1400
rect -906 -1434 -873 -1400
rect -974 -1468 -873 -1434
rect -974 -1502 -940 -1468
rect -906 -1502 -873 -1468
rect -974 -1702 -873 -1502
rect -974 -1736 -940 -1702
rect -906 -1736 -873 -1702
rect -974 -1770 -873 -1736
rect -974 -1804 -940 -1770
rect -906 -1804 -873 -1770
rect -974 -1838 -873 -1804
rect -331 -1400 -230 -1366
rect -331 -1434 -298 -1400
rect -264 -1434 -230 -1400
rect -331 -1468 -230 -1434
rect -331 -1502 -298 -1468
rect -264 -1502 -230 -1468
rect -331 -1702 -230 -1502
rect -331 -1736 -298 -1702
rect -264 -1736 -230 -1702
rect -331 -1770 -230 -1736
rect -331 -1804 -298 -1770
rect -264 -1804 -230 -1770
rect -974 -1872 -940 -1838
rect -906 -1872 -873 -1838
rect -974 -1873 -873 -1872
rect -331 -1838 -230 -1804
rect -331 -1872 -298 -1838
rect -264 -1872 -230 -1838
rect -331 -1873 -230 -1872
rect -974 -1906 -230 -1873
rect -974 -1940 -940 -1906
rect -906 -1940 -872 -1906
rect -838 -1940 -804 -1906
rect -770 -1940 -736 -1906
rect -702 -1940 -502 -1906
rect -468 -1940 -434 -1906
rect -400 -1940 -366 -1906
rect -332 -1940 -298 -1906
rect -264 -1940 -230 -1906
rect -974 -1974 -230 -1940
rect 26 -1264 770 -1230
rect 26 -1298 60 -1264
rect 94 -1298 128 -1264
rect 162 -1298 196 -1264
rect 230 -1298 264 -1264
rect 298 -1298 498 -1264
rect 532 -1298 566 -1264
rect 600 -1298 634 -1264
rect 668 -1298 702 -1264
rect 736 -1298 770 -1264
rect 26 -1331 770 -1298
rect 26 -1332 127 -1331
rect 26 -1366 60 -1332
rect 94 -1366 127 -1332
rect 26 -1400 127 -1366
rect 669 -1332 770 -1331
rect 669 -1366 702 -1332
rect 736 -1366 770 -1332
rect 26 -1434 60 -1400
rect 94 -1434 127 -1400
rect 26 -1468 127 -1434
rect 26 -1502 60 -1468
rect 94 -1502 127 -1468
rect 26 -1702 127 -1502
rect 26 -1736 60 -1702
rect 94 -1736 127 -1702
rect 26 -1770 127 -1736
rect 26 -1804 60 -1770
rect 94 -1804 127 -1770
rect 26 -1838 127 -1804
rect 669 -1400 770 -1366
rect 669 -1434 702 -1400
rect 736 -1434 770 -1400
rect 669 -1468 770 -1434
rect 669 -1502 702 -1468
rect 736 -1502 770 -1468
rect 669 -1702 770 -1502
rect 669 -1736 702 -1702
rect 736 -1736 770 -1702
rect 669 -1770 770 -1736
rect 669 -1804 702 -1770
rect 736 -1804 770 -1770
rect 26 -1872 60 -1838
rect 94 -1872 127 -1838
rect 26 -1873 127 -1872
rect 669 -1838 770 -1804
rect 669 -1872 702 -1838
rect 736 -1872 770 -1838
rect 669 -1873 770 -1872
rect 26 -1906 770 -1873
rect 26 -1940 60 -1906
rect 94 -1940 128 -1906
rect 162 -1940 196 -1906
rect 230 -1940 264 -1906
rect 298 -1940 498 -1906
rect 532 -1940 566 -1906
rect 600 -1940 634 -1906
rect 668 -1940 702 -1906
rect 736 -1940 770 -1906
rect 26 -1974 770 -1940
rect 1026 -1264 1770 -1230
rect 1026 -1298 1060 -1264
rect 1094 -1298 1128 -1264
rect 1162 -1298 1196 -1264
rect 1230 -1298 1264 -1264
rect 1298 -1298 1498 -1264
rect 1532 -1298 1566 -1264
rect 1600 -1298 1634 -1264
rect 1668 -1298 1702 -1264
rect 1736 -1298 1770 -1264
rect 1026 -1331 1770 -1298
rect 1026 -1332 1127 -1331
rect 1026 -1366 1060 -1332
rect 1094 -1366 1127 -1332
rect 1026 -1400 1127 -1366
rect 1669 -1332 1770 -1331
rect 1669 -1366 1702 -1332
rect 1736 -1366 1770 -1332
rect 1026 -1434 1060 -1400
rect 1094 -1434 1127 -1400
rect 1026 -1468 1127 -1434
rect 1026 -1502 1060 -1468
rect 1094 -1502 1127 -1468
rect 1026 -1702 1127 -1502
rect 1026 -1736 1060 -1702
rect 1094 -1736 1127 -1702
rect 1026 -1770 1127 -1736
rect 1026 -1804 1060 -1770
rect 1094 -1804 1127 -1770
rect 1026 -1838 1127 -1804
rect 1669 -1400 1770 -1366
rect 1669 -1434 1702 -1400
rect 1736 -1434 1770 -1400
rect 1669 -1468 1770 -1434
rect 1669 -1502 1702 -1468
rect 1736 -1502 1770 -1468
rect 1669 -1702 1770 -1502
rect 1669 -1736 1702 -1702
rect 1736 -1736 1770 -1702
rect 1669 -1770 1770 -1736
rect 1669 -1804 1702 -1770
rect 1736 -1804 1770 -1770
rect 1026 -1872 1060 -1838
rect 1094 -1872 1127 -1838
rect 1026 -1873 1127 -1872
rect 1669 -1838 1770 -1804
rect 1669 -1872 1702 -1838
rect 1736 -1872 1770 -1838
rect 1669 -1873 1770 -1872
rect 1026 -1906 1770 -1873
rect 1026 -1940 1060 -1906
rect 1094 -1940 1128 -1906
rect 1162 -1940 1196 -1906
rect 1230 -1940 1264 -1906
rect 1298 -1940 1498 -1906
rect 1532 -1940 1566 -1906
rect 1600 -1940 1634 -1906
rect 1668 -1940 1702 -1906
rect 1736 -1940 1770 -1906
rect 1026 -1974 1770 -1940
rect -3974 -2264 -3230 -2230
rect -3974 -2298 -3940 -2264
rect -3906 -2298 -3872 -2264
rect -3838 -2298 -3804 -2264
rect -3770 -2298 -3736 -2264
rect -3702 -2298 -3502 -2264
rect -3468 -2298 -3434 -2264
rect -3400 -2298 -3366 -2264
rect -3332 -2298 -3298 -2264
rect -3264 -2298 -3230 -2264
rect -3974 -2331 -3230 -2298
rect -3974 -2332 -3873 -2331
rect -3974 -2366 -3940 -2332
rect -3906 -2366 -3873 -2332
rect -3974 -2400 -3873 -2366
rect -3331 -2332 -3230 -2331
rect -3331 -2366 -3298 -2332
rect -3264 -2366 -3230 -2332
rect -3974 -2434 -3940 -2400
rect -3906 -2434 -3873 -2400
rect -3974 -2468 -3873 -2434
rect -3974 -2502 -3940 -2468
rect -3906 -2502 -3873 -2468
rect -3974 -2702 -3873 -2502
rect -3974 -2736 -3940 -2702
rect -3906 -2736 -3873 -2702
rect -3974 -2770 -3873 -2736
rect -3974 -2804 -3940 -2770
rect -3906 -2804 -3873 -2770
rect -3974 -2838 -3873 -2804
rect -3331 -2400 -3230 -2366
rect -3331 -2434 -3298 -2400
rect -3264 -2434 -3230 -2400
rect -3331 -2468 -3230 -2434
rect -3331 -2502 -3298 -2468
rect -3264 -2502 -3230 -2468
rect -3331 -2702 -3230 -2502
rect -3331 -2736 -3298 -2702
rect -3264 -2736 -3230 -2702
rect -3331 -2770 -3230 -2736
rect -3331 -2804 -3298 -2770
rect -3264 -2804 -3230 -2770
rect -3974 -2872 -3940 -2838
rect -3906 -2872 -3873 -2838
rect -3974 -2873 -3873 -2872
rect -3331 -2838 -3230 -2804
rect -3331 -2872 -3298 -2838
rect -3264 -2872 -3230 -2838
rect -3331 -2873 -3230 -2872
rect -3974 -2906 -3230 -2873
rect -3974 -2940 -3940 -2906
rect -3906 -2940 -3872 -2906
rect -3838 -2940 -3804 -2906
rect -3770 -2940 -3736 -2906
rect -3702 -2940 -3502 -2906
rect -3468 -2940 -3434 -2906
rect -3400 -2940 -3366 -2906
rect -3332 -2940 -3298 -2906
rect -3264 -2940 -3230 -2906
rect -3974 -2974 -3230 -2940
rect -2974 -2264 -2230 -2230
rect -2974 -2298 -2940 -2264
rect -2906 -2298 -2872 -2264
rect -2838 -2298 -2804 -2264
rect -2770 -2298 -2736 -2264
rect -2702 -2298 -2502 -2264
rect -2468 -2298 -2434 -2264
rect -2400 -2298 -2366 -2264
rect -2332 -2298 -2298 -2264
rect -2264 -2298 -2230 -2264
rect -2974 -2331 -2230 -2298
rect -2974 -2332 -2873 -2331
rect -2974 -2366 -2940 -2332
rect -2906 -2366 -2873 -2332
rect -2974 -2400 -2873 -2366
rect -2331 -2332 -2230 -2331
rect -2331 -2366 -2298 -2332
rect -2264 -2366 -2230 -2332
rect -2974 -2434 -2940 -2400
rect -2906 -2434 -2873 -2400
rect -2974 -2468 -2873 -2434
rect -2974 -2502 -2940 -2468
rect -2906 -2502 -2873 -2468
rect -2974 -2702 -2873 -2502
rect -2974 -2736 -2940 -2702
rect -2906 -2736 -2873 -2702
rect -2974 -2770 -2873 -2736
rect -2974 -2804 -2940 -2770
rect -2906 -2804 -2873 -2770
rect -2974 -2838 -2873 -2804
rect -2331 -2400 -2230 -2366
rect -2331 -2434 -2298 -2400
rect -2264 -2434 -2230 -2400
rect -2331 -2468 -2230 -2434
rect -2331 -2502 -2298 -2468
rect -2264 -2502 -2230 -2468
rect -2331 -2702 -2230 -2502
rect -2331 -2736 -2298 -2702
rect -2264 -2736 -2230 -2702
rect -2331 -2770 -2230 -2736
rect -2331 -2804 -2298 -2770
rect -2264 -2804 -2230 -2770
rect -2974 -2872 -2940 -2838
rect -2906 -2872 -2873 -2838
rect -2974 -2873 -2873 -2872
rect -2331 -2838 -2230 -2804
rect -2331 -2872 -2298 -2838
rect -2264 -2872 -2230 -2838
rect -2331 -2873 -2230 -2872
rect -2974 -2906 -2230 -2873
rect -2974 -2940 -2940 -2906
rect -2906 -2940 -2872 -2906
rect -2838 -2940 -2804 -2906
rect -2770 -2940 -2736 -2906
rect -2702 -2940 -2502 -2906
rect -2468 -2940 -2434 -2906
rect -2400 -2940 -2366 -2906
rect -2332 -2940 -2298 -2906
rect -2264 -2940 -2230 -2906
rect -2974 -2974 -2230 -2940
rect -1974 -2264 -1230 -2230
rect -1974 -2298 -1940 -2264
rect -1906 -2298 -1872 -2264
rect -1838 -2298 -1804 -2264
rect -1770 -2298 -1736 -2264
rect -1702 -2298 -1502 -2264
rect -1468 -2298 -1434 -2264
rect -1400 -2298 -1366 -2264
rect -1332 -2298 -1298 -2264
rect -1264 -2298 -1230 -2264
rect -1974 -2331 -1230 -2298
rect -1974 -2332 -1873 -2331
rect -1974 -2366 -1940 -2332
rect -1906 -2366 -1873 -2332
rect -1974 -2400 -1873 -2366
rect -1331 -2332 -1230 -2331
rect -1331 -2366 -1298 -2332
rect -1264 -2366 -1230 -2332
rect -1974 -2434 -1940 -2400
rect -1906 -2434 -1873 -2400
rect -1974 -2468 -1873 -2434
rect -1974 -2502 -1940 -2468
rect -1906 -2502 -1873 -2468
rect -1974 -2702 -1873 -2502
rect -1974 -2736 -1940 -2702
rect -1906 -2736 -1873 -2702
rect -1974 -2770 -1873 -2736
rect -1974 -2804 -1940 -2770
rect -1906 -2804 -1873 -2770
rect -1974 -2838 -1873 -2804
rect -1331 -2400 -1230 -2366
rect -1331 -2434 -1298 -2400
rect -1264 -2434 -1230 -2400
rect -1331 -2468 -1230 -2434
rect -1331 -2502 -1298 -2468
rect -1264 -2502 -1230 -2468
rect -1331 -2702 -1230 -2502
rect -1331 -2736 -1298 -2702
rect -1264 -2736 -1230 -2702
rect -1331 -2770 -1230 -2736
rect -1331 -2804 -1298 -2770
rect -1264 -2804 -1230 -2770
rect -1974 -2872 -1940 -2838
rect -1906 -2872 -1873 -2838
rect -1974 -2873 -1873 -2872
rect -1331 -2838 -1230 -2804
rect -1331 -2872 -1298 -2838
rect -1264 -2872 -1230 -2838
rect -1331 -2873 -1230 -2872
rect -1974 -2906 -1230 -2873
rect -1974 -2940 -1940 -2906
rect -1906 -2940 -1872 -2906
rect -1838 -2940 -1804 -2906
rect -1770 -2940 -1736 -2906
rect -1702 -2940 -1502 -2906
rect -1468 -2940 -1434 -2906
rect -1400 -2940 -1366 -2906
rect -1332 -2940 -1298 -2906
rect -1264 -2940 -1230 -2906
rect -1974 -2974 -1230 -2940
rect -974 -2264 -230 -2230
rect -974 -2298 -940 -2264
rect -906 -2298 -872 -2264
rect -838 -2298 -804 -2264
rect -770 -2298 -736 -2264
rect -702 -2298 -502 -2264
rect -468 -2298 -434 -2264
rect -400 -2298 -366 -2264
rect -332 -2298 -298 -2264
rect -264 -2298 -230 -2264
rect -974 -2331 -230 -2298
rect -974 -2332 -873 -2331
rect -974 -2366 -940 -2332
rect -906 -2366 -873 -2332
rect -974 -2400 -873 -2366
rect -331 -2332 -230 -2331
rect -331 -2366 -298 -2332
rect -264 -2366 -230 -2332
rect -974 -2434 -940 -2400
rect -906 -2434 -873 -2400
rect -974 -2468 -873 -2434
rect -974 -2502 -940 -2468
rect -906 -2502 -873 -2468
rect -974 -2702 -873 -2502
rect -974 -2736 -940 -2702
rect -906 -2736 -873 -2702
rect -974 -2770 -873 -2736
rect -974 -2804 -940 -2770
rect -906 -2804 -873 -2770
rect -974 -2838 -873 -2804
rect -331 -2400 -230 -2366
rect -331 -2434 -298 -2400
rect -264 -2434 -230 -2400
rect -331 -2468 -230 -2434
rect -331 -2502 -298 -2468
rect -264 -2502 -230 -2468
rect -331 -2702 -230 -2502
rect -331 -2736 -298 -2702
rect -264 -2736 -230 -2702
rect -331 -2770 -230 -2736
rect -331 -2804 -298 -2770
rect -264 -2804 -230 -2770
rect -974 -2872 -940 -2838
rect -906 -2872 -873 -2838
rect -974 -2873 -873 -2872
rect -331 -2838 -230 -2804
rect -331 -2872 -298 -2838
rect -264 -2872 -230 -2838
rect -331 -2873 -230 -2872
rect -974 -2906 -230 -2873
rect -974 -2940 -940 -2906
rect -906 -2940 -872 -2906
rect -838 -2940 -804 -2906
rect -770 -2940 -736 -2906
rect -702 -2940 -502 -2906
rect -468 -2940 -434 -2906
rect -400 -2940 -366 -2906
rect -332 -2940 -298 -2906
rect -264 -2940 -230 -2906
rect -974 -2974 -230 -2940
rect 26 -2264 770 -2230
rect 26 -2298 60 -2264
rect 94 -2298 128 -2264
rect 162 -2298 196 -2264
rect 230 -2298 264 -2264
rect 298 -2298 498 -2264
rect 532 -2298 566 -2264
rect 600 -2298 634 -2264
rect 668 -2298 702 -2264
rect 736 -2298 770 -2264
rect 26 -2331 770 -2298
rect 26 -2332 127 -2331
rect 26 -2366 60 -2332
rect 94 -2366 127 -2332
rect 26 -2400 127 -2366
rect 669 -2332 770 -2331
rect 669 -2366 702 -2332
rect 736 -2366 770 -2332
rect 26 -2434 60 -2400
rect 94 -2434 127 -2400
rect 26 -2468 127 -2434
rect 26 -2502 60 -2468
rect 94 -2502 127 -2468
rect 26 -2702 127 -2502
rect 26 -2736 60 -2702
rect 94 -2736 127 -2702
rect 26 -2770 127 -2736
rect 26 -2804 60 -2770
rect 94 -2804 127 -2770
rect 26 -2838 127 -2804
rect 669 -2400 770 -2366
rect 669 -2434 702 -2400
rect 736 -2434 770 -2400
rect 669 -2468 770 -2434
rect 669 -2502 702 -2468
rect 736 -2502 770 -2468
rect 669 -2702 770 -2502
rect 669 -2736 702 -2702
rect 736 -2736 770 -2702
rect 669 -2770 770 -2736
rect 669 -2804 702 -2770
rect 736 -2804 770 -2770
rect 26 -2872 60 -2838
rect 94 -2872 127 -2838
rect 26 -2873 127 -2872
rect 669 -2838 770 -2804
rect 669 -2872 702 -2838
rect 736 -2872 770 -2838
rect 669 -2873 770 -2872
rect 26 -2906 770 -2873
rect 26 -2940 60 -2906
rect 94 -2940 128 -2906
rect 162 -2940 196 -2906
rect 230 -2940 264 -2906
rect 298 -2940 498 -2906
rect 532 -2940 566 -2906
rect 600 -2940 634 -2906
rect 668 -2940 702 -2906
rect 736 -2940 770 -2906
rect 26 -2974 770 -2940
rect 1026 -2264 1770 -2230
rect 1026 -2298 1060 -2264
rect 1094 -2298 1128 -2264
rect 1162 -2298 1196 -2264
rect 1230 -2298 1264 -2264
rect 1298 -2298 1498 -2264
rect 1532 -2298 1566 -2264
rect 1600 -2298 1634 -2264
rect 1668 -2298 1702 -2264
rect 1736 -2298 1770 -2264
rect 1026 -2331 1770 -2298
rect 1026 -2332 1127 -2331
rect 1026 -2366 1060 -2332
rect 1094 -2366 1127 -2332
rect 1026 -2400 1127 -2366
rect 1669 -2332 1770 -2331
rect 1669 -2366 1702 -2332
rect 1736 -2366 1770 -2332
rect 1026 -2434 1060 -2400
rect 1094 -2434 1127 -2400
rect 1026 -2468 1127 -2434
rect 1026 -2502 1060 -2468
rect 1094 -2502 1127 -2468
rect 1026 -2702 1127 -2502
rect 1026 -2736 1060 -2702
rect 1094 -2736 1127 -2702
rect 1026 -2770 1127 -2736
rect 1026 -2804 1060 -2770
rect 1094 -2804 1127 -2770
rect 1026 -2838 1127 -2804
rect 1669 -2400 1770 -2366
rect 1669 -2434 1702 -2400
rect 1736 -2434 1770 -2400
rect 1669 -2468 1770 -2434
rect 1669 -2502 1702 -2468
rect 1736 -2502 1770 -2468
rect 1669 -2702 1770 -2502
rect 1669 -2736 1702 -2702
rect 1736 -2736 1770 -2702
rect 1669 -2770 1770 -2736
rect 1669 -2804 1702 -2770
rect 1736 -2804 1770 -2770
rect 1026 -2872 1060 -2838
rect 1094 -2872 1127 -2838
rect 1026 -2873 1127 -2872
rect 1669 -2838 1770 -2804
rect 1669 -2872 1702 -2838
rect 1736 -2872 1770 -2838
rect 1669 -2873 1770 -2872
rect 1026 -2906 1770 -2873
rect 1026 -2940 1060 -2906
rect 1094 -2940 1128 -2906
rect 1162 -2940 1196 -2906
rect 1230 -2940 1264 -2906
rect 1298 -2940 1498 -2906
rect 1532 -2940 1566 -2906
rect 1600 -2940 1634 -2906
rect 1668 -2940 1702 -2906
rect 1736 -2940 1770 -2906
rect 1026 -2974 1770 -2940
<< nsubdiff >>
rect -3811 1583 -3393 1607
rect -3811 1549 -3787 1583
rect -3753 1549 -3719 1583
rect -3685 1549 -3519 1583
rect -3485 1549 -3451 1583
rect -3417 1549 -3393 1583
rect -3811 1535 -3393 1549
rect -3811 1515 -3739 1535
rect -3811 1481 -3787 1515
rect -3753 1481 -3739 1515
rect -3811 1315 -3739 1481
rect -3465 1515 -3393 1535
rect -3465 1481 -3451 1515
rect -3417 1481 -3393 1515
rect -3811 1281 -3787 1315
rect -3753 1281 -3739 1315
rect -3811 1261 -3739 1281
rect -3465 1315 -3393 1481
rect -3465 1281 -3451 1315
rect -3417 1281 -3393 1315
rect -3465 1261 -3393 1281
rect -3811 1247 -3393 1261
rect -3811 1213 -3787 1247
rect -3753 1213 -3719 1247
rect -3685 1213 -3519 1247
rect -3485 1213 -3451 1247
rect -3417 1213 -3393 1247
rect -3811 1189 -3393 1213
rect -2811 1583 -2393 1607
rect -2811 1549 -2787 1583
rect -2753 1549 -2719 1583
rect -2685 1549 -2519 1583
rect -2485 1549 -2451 1583
rect -2417 1549 -2393 1583
rect -2811 1535 -2393 1549
rect -2811 1515 -2739 1535
rect -2811 1481 -2787 1515
rect -2753 1481 -2739 1515
rect -2811 1315 -2739 1481
rect -2465 1515 -2393 1535
rect -2465 1481 -2451 1515
rect -2417 1481 -2393 1515
rect -2811 1281 -2787 1315
rect -2753 1281 -2739 1315
rect -2811 1261 -2739 1281
rect -2465 1315 -2393 1481
rect -2465 1281 -2451 1315
rect -2417 1281 -2393 1315
rect -2465 1261 -2393 1281
rect -2811 1247 -2393 1261
rect -2811 1213 -2787 1247
rect -2753 1213 -2719 1247
rect -2685 1213 -2519 1247
rect -2485 1213 -2451 1247
rect -2417 1213 -2393 1247
rect -2811 1189 -2393 1213
rect -1811 1583 -1393 1607
rect -1811 1549 -1787 1583
rect -1753 1549 -1719 1583
rect -1685 1549 -1519 1583
rect -1485 1549 -1451 1583
rect -1417 1549 -1393 1583
rect -1811 1535 -1393 1549
rect -1811 1515 -1739 1535
rect -1811 1481 -1787 1515
rect -1753 1481 -1739 1515
rect -1811 1315 -1739 1481
rect -1465 1515 -1393 1535
rect -1465 1481 -1451 1515
rect -1417 1481 -1393 1515
rect -1811 1281 -1787 1315
rect -1753 1281 -1739 1315
rect -1811 1261 -1739 1281
rect -1465 1315 -1393 1481
rect -1465 1281 -1451 1315
rect -1417 1281 -1393 1315
rect -1465 1261 -1393 1281
rect -1811 1247 -1393 1261
rect -1811 1213 -1787 1247
rect -1753 1213 -1719 1247
rect -1685 1213 -1519 1247
rect -1485 1213 -1451 1247
rect -1417 1213 -1393 1247
rect -1811 1189 -1393 1213
rect -811 1583 -393 1607
rect -811 1549 -787 1583
rect -753 1549 -719 1583
rect -685 1549 -519 1583
rect -485 1549 -451 1583
rect -417 1549 -393 1583
rect -811 1535 -393 1549
rect -811 1515 -739 1535
rect -811 1481 -787 1515
rect -753 1481 -739 1515
rect -811 1315 -739 1481
rect -465 1515 -393 1535
rect -465 1481 -451 1515
rect -417 1481 -393 1515
rect -811 1281 -787 1315
rect -753 1281 -739 1315
rect -811 1261 -739 1281
rect -465 1315 -393 1481
rect -465 1281 -451 1315
rect -417 1281 -393 1315
rect -465 1261 -393 1281
rect -811 1247 -393 1261
rect -811 1213 -787 1247
rect -753 1213 -719 1247
rect -685 1213 -519 1247
rect -485 1213 -451 1247
rect -417 1213 -393 1247
rect -811 1189 -393 1213
rect 189 1583 607 1607
rect 189 1549 213 1583
rect 247 1549 281 1583
rect 315 1549 481 1583
rect 515 1549 549 1583
rect 583 1549 607 1583
rect 189 1535 607 1549
rect 189 1515 261 1535
rect 189 1481 213 1515
rect 247 1481 261 1515
rect 189 1315 261 1481
rect 535 1515 607 1535
rect 535 1481 549 1515
rect 583 1481 607 1515
rect 189 1281 213 1315
rect 247 1281 261 1315
rect 189 1261 261 1281
rect 535 1315 607 1481
rect 535 1281 549 1315
rect 583 1281 607 1315
rect 535 1261 607 1281
rect 189 1247 607 1261
rect 189 1213 213 1247
rect 247 1213 281 1247
rect 315 1213 481 1247
rect 515 1213 549 1247
rect 583 1213 607 1247
rect 189 1189 607 1213
rect 1189 1583 1607 1607
rect 1189 1549 1213 1583
rect 1247 1549 1281 1583
rect 1315 1549 1481 1583
rect 1515 1549 1549 1583
rect 1583 1549 1607 1583
rect 1189 1535 1607 1549
rect 1189 1515 1261 1535
rect 1189 1481 1213 1515
rect 1247 1481 1261 1515
rect 1189 1315 1261 1481
rect 1535 1515 1607 1535
rect 1535 1481 1549 1515
rect 1583 1481 1607 1515
rect 1189 1281 1213 1315
rect 1247 1281 1261 1315
rect 1189 1261 1261 1281
rect 1535 1315 1607 1481
rect 1535 1281 1549 1315
rect 1583 1281 1607 1315
rect 1535 1261 1607 1281
rect 1189 1247 1607 1261
rect 1189 1213 1213 1247
rect 1247 1213 1281 1247
rect 1315 1213 1481 1247
rect 1515 1213 1549 1247
rect 1583 1213 1607 1247
rect 1189 1189 1607 1213
rect -3811 583 -3393 607
rect -3811 549 -3787 583
rect -3753 549 -3719 583
rect -3685 549 -3519 583
rect -3485 549 -3451 583
rect -3417 549 -3393 583
rect -3811 535 -3393 549
rect -3811 515 -3739 535
rect -3811 481 -3787 515
rect -3753 481 -3739 515
rect -3811 315 -3739 481
rect -3465 515 -3393 535
rect -3465 481 -3451 515
rect -3417 481 -3393 515
rect -3811 281 -3787 315
rect -3753 281 -3739 315
rect -3811 261 -3739 281
rect -3465 315 -3393 481
rect -3465 281 -3451 315
rect -3417 281 -3393 315
rect -3465 261 -3393 281
rect -3811 247 -3393 261
rect -3811 213 -3787 247
rect -3753 213 -3719 247
rect -3685 213 -3519 247
rect -3485 213 -3451 247
rect -3417 213 -3393 247
rect -3811 189 -3393 213
rect -2811 583 -2393 607
rect -2811 549 -2787 583
rect -2753 549 -2719 583
rect -2685 549 -2519 583
rect -2485 549 -2451 583
rect -2417 549 -2393 583
rect -2811 535 -2393 549
rect -2811 515 -2739 535
rect -2811 481 -2787 515
rect -2753 481 -2739 515
rect -2811 315 -2739 481
rect -2465 515 -2393 535
rect -2465 481 -2451 515
rect -2417 481 -2393 515
rect -2811 281 -2787 315
rect -2753 281 -2739 315
rect -2811 261 -2739 281
rect -2465 315 -2393 481
rect -2465 281 -2451 315
rect -2417 281 -2393 315
rect -2465 261 -2393 281
rect -2811 247 -2393 261
rect -2811 213 -2787 247
rect -2753 213 -2719 247
rect -2685 213 -2519 247
rect -2485 213 -2451 247
rect -2417 213 -2393 247
rect -2811 189 -2393 213
rect -1811 583 -1393 607
rect -1811 549 -1787 583
rect -1753 549 -1719 583
rect -1685 549 -1519 583
rect -1485 549 -1451 583
rect -1417 549 -1393 583
rect -1811 535 -1393 549
rect -1811 515 -1739 535
rect -1811 481 -1787 515
rect -1753 481 -1739 515
rect -1811 315 -1739 481
rect -1465 515 -1393 535
rect -1465 481 -1451 515
rect -1417 481 -1393 515
rect -1811 281 -1787 315
rect -1753 281 -1739 315
rect -1811 261 -1739 281
rect -1465 315 -1393 481
rect -1465 281 -1451 315
rect -1417 281 -1393 315
rect -1465 261 -1393 281
rect -1811 247 -1393 261
rect -1811 213 -1787 247
rect -1753 213 -1719 247
rect -1685 213 -1519 247
rect -1485 213 -1451 247
rect -1417 213 -1393 247
rect -1811 189 -1393 213
rect -811 583 -393 607
rect -811 549 -787 583
rect -753 549 -719 583
rect -685 549 -519 583
rect -485 549 -451 583
rect -417 549 -393 583
rect -811 535 -393 549
rect -811 515 -739 535
rect -811 481 -787 515
rect -753 481 -739 515
rect -811 315 -739 481
rect -465 515 -393 535
rect -465 481 -451 515
rect -417 481 -393 515
rect -811 281 -787 315
rect -753 281 -739 315
rect -811 261 -739 281
rect -465 315 -393 481
rect -465 281 -451 315
rect -417 281 -393 315
rect -465 261 -393 281
rect -811 247 -393 261
rect -811 213 -787 247
rect -753 213 -719 247
rect -685 213 -519 247
rect -485 213 -451 247
rect -417 213 -393 247
rect -811 189 -393 213
rect 189 583 607 607
rect 189 549 213 583
rect 247 549 281 583
rect 315 549 481 583
rect 515 549 549 583
rect 583 549 607 583
rect 189 535 607 549
rect 189 515 261 535
rect 189 481 213 515
rect 247 481 261 515
rect 189 315 261 481
rect 535 515 607 535
rect 535 481 549 515
rect 583 481 607 515
rect 189 281 213 315
rect 247 281 261 315
rect 189 261 261 281
rect 535 315 607 481
rect 535 281 549 315
rect 583 281 607 315
rect 535 261 607 281
rect 189 247 607 261
rect 189 213 213 247
rect 247 213 281 247
rect 315 213 481 247
rect 515 213 549 247
rect 583 213 607 247
rect 189 189 607 213
rect 1189 583 1607 607
rect 1189 549 1213 583
rect 1247 549 1281 583
rect 1315 549 1481 583
rect 1515 549 1549 583
rect 1583 549 1607 583
rect 1189 535 1607 549
rect 1189 515 1261 535
rect 1189 481 1213 515
rect 1247 481 1261 515
rect 1189 315 1261 481
rect 1535 515 1607 535
rect 1535 481 1549 515
rect 1583 481 1607 515
rect 1189 281 1213 315
rect 1247 281 1261 315
rect 1189 261 1261 281
rect 1535 315 1607 481
rect 1535 281 1549 315
rect 1583 281 1607 315
rect 1535 261 1607 281
rect 1189 247 1607 261
rect 1189 213 1213 247
rect 1247 213 1281 247
rect 1315 213 1481 247
rect 1515 213 1549 247
rect 1583 213 1607 247
rect 1189 189 1607 213
rect -3811 -417 -3393 -393
rect -3811 -451 -3787 -417
rect -3753 -451 -3719 -417
rect -3685 -451 -3519 -417
rect -3485 -451 -3451 -417
rect -3417 -451 -3393 -417
rect -3811 -465 -3393 -451
rect -3811 -485 -3739 -465
rect -3811 -519 -3787 -485
rect -3753 -519 -3739 -485
rect -3811 -685 -3739 -519
rect -3465 -485 -3393 -465
rect -3465 -519 -3451 -485
rect -3417 -519 -3393 -485
rect -3811 -719 -3787 -685
rect -3753 -719 -3739 -685
rect -3811 -739 -3739 -719
rect -3465 -685 -3393 -519
rect -3465 -719 -3451 -685
rect -3417 -719 -3393 -685
rect -3465 -739 -3393 -719
rect -3811 -753 -3393 -739
rect -3811 -787 -3787 -753
rect -3753 -787 -3719 -753
rect -3685 -787 -3519 -753
rect -3485 -787 -3451 -753
rect -3417 -787 -3393 -753
rect -3811 -811 -3393 -787
rect -2811 -417 -2393 -393
rect -2811 -451 -2787 -417
rect -2753 -451 -2719 -417
rect -2685 -451 -2519 -417
rect -2485 -451 -2451 -417
rect -2417 -451 -2393 -417
rect -2811 -465 -2393 -451
rect -2811 -485 -2739 -465
rect -2811 -519 -2787 -485
rect -2753 -519 -2739 -485
rect -2811 -685 -2739 -519
rect -2465 -485 -2393 -465
rect -2465 -519 -2451 -485
rect -2417 -519 -2393 -485
rect -2811 -719 -2787 -685
rect -2753 -719 -2739 -685
rect -2811 -739 -2739 -719
rect -2465 -685 -2393 -519
rect -2465 -719 -2451 -685
rect -2417 -719 -2393 -685
rect -2465 -739 -2393 -719
rect -2811 -753 -2393 -739
rect -2811 -787 -2787 -753
rect -2753 -787 -2719 -753
rect -2685 -787 -2519 -753
rect -2485 -787 -2451 -753
rect -2417 -787 -2393 -753
rect -2811 -811 -2393 -787
rect -1811 -417 -1393 -393
rect -1811 -451 -1787 -417
rect -1753 -451 -1719 -417
rect -1685 -451 -1519 -417
rect -1485 -451 -1451 -417
rect -1417 -451 -1393 -417
rect -1811 -465 -1393 -451
rect -1811 -485 -1739 -465
rect -1811 -519 -1787 -485
rect -1753 -519 -1739 -485
rect -1811 -685 -1739 -519
rect -1465 -485 -1393 -465
rect -1465 -519 -1451 -485
rect -1417 -519 -1393 -485
rect -1811 -719 -1787 -685
rect -1753 -719 -1739 -685
rect -1811 -739 -1739 -719
rect -1465 -685 -1393 -519
rect -1465 -719 -1451 -685
rect -1417 -719 -1393 -685
rect -1465 -739 -1393 -719
rect -1811 -753 -1393 -739
rect -1811 -787 -1787 -753
rect -1753 -787 -1719 -753
rect -1685 -787 -1519 -753
rect -1485 -787 -1451 -753
rect -1417 -787 -1393 -753
rect -1811 -811 -1393 -787
rect -811 -417 -393 -393
rect -811 -451 -787 -417
rect -753 -451 -719 -417
rect -685 -451 -519 -417
rect -485 -451 -451 -417
rect -417 -451 -393 -417
rect -811 -465 -393 -451
rect -811 -485 -739 -465
rect -811 -519 -787 -485
rect -753 -519 -739 -485
rect -811 -685 -739 -519
rect -465 -485 -393 -465
rect -465 -519 -451 -485
rect -417 -519 -393 -485
rect -811 -719 -787 -685
rect -753 -719 -739 -685
rect -811 -739 -739 -719
rect -465 -685 -393 -519
rect -465 -719 -451 -685
rect -417 -719 -393 -685
rect -465 -739 -393 -719
rect -811 -753 -393 -739
rect -811 -787 -787 -753
rect -753 -787 -719 -753
rect -685 -787 -519 -753
rect -485 -787 -451 -753
rect -417 -787 -393 -753
rect -811 -811 -393 -787
rect 189 -417 607 -393
rect 189 -451 213 -417
rect 247 -451 281 -417
rect 315 -451 481 -417
rect 515 -451 549 -417
rect 583 -451 607 -417
rect 189 -465 607 -451
rect 189 -485 261 -465
rect 189 -519 213 -485
rect 247 -519 261 -485
rect 189 -685 261 -519
rect 535 -485 607 -465
rect 535 -519 549 -485
rect 583 -519 607 -485
rect 189 -719 213 -685
rect 247 -719 261 -685
rect 189 -739 261 -719
rect 535 -685 607 -519
rect 535 -719 549 -685
rect 583 -719 607 -685
rect 535 -739 607 -719
rect 189 -753 607 -739
rect 189 -787 213 -753
rect 247 -787 281 -753
rect 315 -787 481 -753
rect 515 -787 549 -753
rect 583 -787 607 -753
rect 189 -811 607 -787
rect 1189 -417 1607 -393
rect 1189 -451 1213 -417
rect 1247 -451 1281 -417
rect 1315 -451 1481 -417
rect 1515 -451 1549 -417
rect 1583 -451 1607 -417
rect 1189 -465 1607 -451
rect 1189 -485 1261 -465
rect 1189 -519 1213 -485
rect 1247 -519 1261 -485
rect 1189 -685 1261 -519
rect 1535 -485 1607 -465
rect 1535 -519 1549 -485
rect 1583 -519 1607 -485
rect 1189 -719 1213 -685
rect 1247 -719 1261 -685
rect 1189 -739 1261 -719
rect 1535 -685 1607 -519
rect 1535 -719 1549 -685
rect 1583 -719 1607 -685
rect 1535 -739 1607 -719
rect 1189 -753 1607 -739
rect 1189 -787 1213 -753
rect 1247 -787 1281 -753
rect 1315 -787 1481 -753
rect 1515 -787 1549 -753
rect 1583 -787 1607 -753
rect 1189 -811 1607 -787
rect -3811 -1417 -3393 -1393
rect -3811 -1451 -3787 -1417
rect -3753 -1451 -3719 -1417
rect -3685 -1451 -3519 -1417
rect -3485 -1451 -3451 -1417
rect -3417 -1451 -3393 -1417
rect -3811 -1465 -3393 -1451
rect -3811 -1485 -3739 -1465
rect -3811 -1519 -3787 -1485
rect -3753 -1519 -3739 -1485
rect -3811 -1685 -3739 -1519
rect -3465 -1485 -3393 -1465
rect -3465 -1519 -3451 -1485
rect -3417 -1519 -3393 -1485
rect -3811 -1719 -3787 -1685
rect -3753 -1719 -3739 -1685
rect -3811 -1739 -3739 -1719
rect -3465 -1685 -3393 -1519
rect -3465 -1719 -3451 -1685
rect -3417 -1719 -3393 -1685
rect -3465 -1739 -3393 -1719
rect -3811 -1753 -3393 -1739
rect -3811 -1787 -3787 -1753
rect -3753 -1787 -3719 -1753
rect -3685 -1787 -3519 -1753
rect -3485 -1787 -3451 -1753
rect -3417 -1787 -3393 -1753
rect -3811 -1811 -3393 -1787
rect -2811 -1417 -2393 -1393
rect -2811 -1451 -2787 -1417
rect -2753 -1451 -2719 -1417
rect -2685 -1451 -2519 -1417
rect -2485 -1451 -2451 -1417
rect -2417 -1451 -2393 -1417
rect -2811 -1465 -2393 -1451
rect -2811 -1485 -2739 -1465
rect -2811 -1519 -2787 -1485
rect -2753 -1519 -2739 -1485
rect -2811 -1685 -2739 -1519
rect -2465 -1485 -2393 -1465
rect -2465 -1519 -2451 -1485
rect -2417 -1519 -2393 -1485
rect -2811 -1719 -2787 -1685
rect -2753 -1719 -2739 -1685
rect -2811 -1739 -2739 -1719
rect -2465 -1685 -2393 -1519
rect -2465 -1719 -2451 -1685
rect -2417 -1719 -2393 -1685
rect -2465 -1739 -2393 -1719
rect -2811 -1753 -2393 -1739
rect -2811 -1787 -2787 -1753
rect -2753 -1787 -2719 -1753
rect -2685 -1787 -2519 -1753
rect -2485 -1787 -2451 -1753
rect -2417 -1787 -2393 -1753
rect -2811 -1811 -2393 -1787
rect -1811 -1417 -1393 -1393
rect -1811 -1451 -1787 -1417
rect -1753 -1451 -1719 -1417
rect -1685 -1451 -1519 -1417
rect -1485 -1451 -1451 -1417
rect -1417 -1451 -1393 -1417
rect -1811 -1465 -1393 -1451
rect -1811 -1485 -1739 -1465
rect -1811 -1519 -1787 -1485
rect -1753 -1519 -1739 -1485
rect -1811 -1685 -1739 -1519
rect -1465 -1485 -1393 -1465
rect -1465 -1519 -1451 -1485
rect -1417 -1519 -1393 -1485
rect -1811 -1719 -1787 -1685
rect -1753 -1719 -1739 -1685
rect -1811 -1739 -1739 -1719
rect -1465 -1685 -1393 -1519
rect -1465 -1719 -1451 -1685
rect -1417 -1719 -1393 -1685
rect -1465 -1739 -1393 -1719
rect -1811 -1753 -1393 -1739
rect -1811 -1787 -1787 -1753
rect -1753 -1787 -1719 -1753
rect -1685 -1787 -1519 -1753
rect -1485 -1787 -1451 -1753
rect -1417 -1787 -1393 -1753
rect -1811 -1811 -1393 -1787
rect -811 -1417 -393 -1393
rect -811 -1451 -787 -1417
rect -753 -1451 -719 -1417
rect -685 -1451 -519 -1417
rect -485 -1451 -451 -1417
rect -417 -1451 -393 -1417
rect -811 -1465 -393 -1451
rect -811 -1485 -739 -1465
rect -811 -1519 -787 -1485
rect -753 -1519 -739 -1485
rect -811 -1685 -739 -1519
rect -465 -1485 -393 -1465
rect -465 -1519 -451 -1485
rect -417 -1519 -393 -1485
rect -811 -1719 -787 -1685
rect -753 -1719 -739 -1685
rect -811 -1739 -739 -1719
rect -465 -1685 -393 -1519
rect -465 -1719 -451 -1685
rect -417 -1719 -393 -1685
rect -465 -1739 -393 -1719
rect -811 -1753 -393 -1739
rect -811 -1787 -787 -1753
rect -753 -1787 -719 -1753
rect -685 -1787 -519 -1753
rect -485 -1787 -451 -1753
rect -417 -1787 -393 -1753
rect -811 -1811 -393 -1787
rect 189 -1417 607 -1393
rect 189 -1451 213 -1417
rect 247 -1451 281 -1417
rect 315 -1451 481 -1417
rect 515 -1451 549 -1417
rect 583 -1451 607 -1417
rect 189 -1465 607 -1451
rect 189 -1485 261 -1465
rect 189 -1519 213 -1485
rect 247 -1519 261 -1485
rect 189 -1685 261 -1519
rect 535 -1485 607 -1465
rect 535 -1519 549 -1485
rect 583 -1519 607 -1485
rect 189 -1719 213 -1685
rect 247 -1719 261 -1685
rect 189 -1739 261 -1719
rect 535 -1685 607 -1519
rect 535 -1719 549 -1685
rect 583 -1719 607 -1685
rect 535 -1739 607 -1719
rect 189 -1753 607 -1739
rect 189 -1787 213 -1753
rect 247 -1787 281 -1753
rect 315 -1787 481 -1753
rect 515 -1787 549 -1753
rect 583 -1787 607 -1753
rect 189 -1811 607 -1787
rect 1189 -1417 1607 -1393
rect 1189 -1451 1213 -1417
rect 1247 -1451 1281 -1417
rect 1315 -1451 1481 -1417
rect 1515 -1451 1549 -1417
rect 1583 -1451 1607 -1417
rect 1189 -1465 1607 -1451
rect 1189 -1485 1261 -1465
rect 1189 -1519 1213 -1485
rect 1247 -1519 1261 -1485
rect 1189 -1685 1261 -1519
rect 1535 -1485 1607 -1465
rect 1535 -1519 1549 -1485
rect 1583 -1519 1607 -1485
rect 1189 -1719 1213 -1685
rect 1247 -1719 1261 -1685
rect 1189 -1739 1261 -1719
rect 1535 -1685 1607 -1519
rect 1535 -1719 1549 -1685
rect 1583 -1719 1607 -1685
rect 1535 -1739 1607 -1719
rect 1189 -1753 1607 -1739
rect 1189 -1787 1213 -1753
rect 1247 -1787 1281 -1753
rect 1315 -1787 1481 -1753
rect 1515 -1787 1549 -1753
rect 1583 -1787 1607 -1753
rect 1189 -1811 1607 -1787
rect -3811 -2417 -3393 -2393
rect -3811 -2451 -3787 -2417
rect -3753 -2451 -3719 -2417
rect -3685 -2451 -3519 -2417
rect -3485 -2451 -3451 -2417
rect -3417 -2451 -3393 -2417
rect -3811 -2465 -3393 -2451
rect -3811 -2485 -3739 -2465
rect -3811 -2519 -3787 -2485
rect -3753 -2519 -3739 -2485
rect -3811 -2685 -3739 -2519
rect -3465 -2485 -3393 -2465
rect -3465 -2519 -3451 -2485
rect -3417 -2519 -3393 -2485
rect -3811 -2719 -3787 -2685
rect -3753 -2719 -3739 -2685
rect -3811 -2739 -3739 -2719
rect -3465 -2685 -3393 -2519
rect -3465 -2719 -3451 -2685
rect -3417 -2719 -3393 -2685
rect -3465 -2739 -3393 -2719
rect -3811 -2753 -3393 -2739
rect -3811 -2787 -3787 -2753
rect -3753 -2787 -3719 -2753
rect -3685 -2787 -3519 -2753
rect -3485 -2787 -3451 -2753
rect -3417 -2787 -3393 -2753
rect -3811 -2811 -3393 -2787
rect -2811 -2417 -2393 -2393
rect -2811 -2451 -2787 -2417
rect -2753 -2451 -2719 -2417
rect -2685 -2451 -2519 -2417
rect -2485 -2451 -2451 -2417
rect -2417 -2451 -2393 -2417
rect -2811 -2465 -2393 -2451
rect -2811 -2485 -2739 -2465
rect -2811 -2519 -2787 -2485
rect -2753 -2519 -2739 -2485
rect -2811 -2685 -2739 -2519
rect -2465 -2485 -2393 -2465
rect -2465 -2519 -2451 -2485
rect -2417 -2519 -2393 -2485
rect -2811 -2719 -2787 -2685
rect -2753 -2719 -2739 -2685
rect -2811 -2739 -2739 -2719
rect -2465 -2685 -2393 -2519
rect -2465 -2719 -2451 -2685
rect -2417 -2719 -2393 -2685
rect -2465 -2739 -2393 -2719
rect -2811 -2753 -2393 -2739
rect -2811 -2787 -2787 -2753
rect -2753 -2787 -2719 -2753
rect -2685 -2787 -2519 -2753
rect -2485 -2787 -2451 -2753
rect -2417 -2787 -2393 -2753
rect -2811 -2811 -2393 -2787
rect -1811 -2417 -1393 -2393
rect -1811 -2451 -1787 -2417
rect -1753 -2451 -1719 -2417
rect -1685 -2451 -1519 -2417
rect -1485 -2451 -1451 -2417
rect -1417 -2451 -1393 -2417
rect -1811 -2465 -1393 -2451
rect -1811 -2485 -1739 -2465
rect -1811 -2519 -1787 -2485
rect -1753 -2519 -1739 -2485
rect -1811 -2685 -1739 -2519
rect -1465 -2485 -1393 -2465
rect -1465 -2519 -1451 -2485
rect -1417 -2519 -1393 -2485
rect -1811 -2719 -1787 -2685
rect -1753 -2719 -1739 -2685
rect -1811 -2739 -1739 -2719
rect -1465 -2685 -1393 -2519
rect -1465 -2719 -1451 -2685
rect -1417 -2719 -1393 -2685
rect -1465 -2739 -1393 -2719
rect -1811 -2753 -1393 -2739
rect -1811 -2787 -1787 -2753
rect -1753 -2787 -1719 -2753
rect -1685 -2787 -1519 -2753
rect -1485 -2787 -1451 -2753
rect -1417 -2787 -1393 -2753
rect -1811 -2811 -1393 -2787
rect -811 -2417 -393 -2393
rect -811 -2451 -787 -2417
rect -753 -2451 -719 -2417
rect -685 -2451 -519 -2417
rect -485 -2451 -451 -2417
rect -417 -2451 -393 -2417
rect -811 -2465 -393 -2451
rect -811 -2485 -739 -2465
rect -811 -2519 -787 -2485
rect -753 -2519 -739 -2485
rect -811 -2685 -739 -2519
rect -465 -2485 -393 -2465
rect -465 -2519 -451 -2485
rect -417 -2519 -393 -2485
rect -811 -2719 -787 -2685
rect -753 -2719 -739 -2685
rect -811 -2739 -739 -2719
rect -465 -2685 -393 -2519
rect -465 -2719 -451 -2685
rect -417 -2719 -393 -2685
rect -465 -2739 -393 -2719
rect -811 -2753 -393 -2739
rect -811 -2787 -787 -2753
rect -753 -2787 -719 -2753
rect -685 -2787 -519 -2753
rect -485 -2787 -451 -2753
rect -417 -2787 -393 -2753
rect -811 -2811 -393 -2787
rect 189 -2417 607 -2393
rect 189 -2451 213 -2417
rect 247 -2451 281 -2417
rect 315 -2451 481 -2417
rect 515 -2451 549 -2417
rect 583 -2451 607 -2417
rect 189 -2465 607 -2451
rect 189 -2485 261 -2465
rect 189 -2519 213 -2485
rect 247 -2519 261 -2485
rect 189 -2685 261 -2519
rect 535 -2485 607 -2465
rect 535 -2519 549 -2485
rect 583 -2519 607 -2485
rect 189 -2719 213 -2685
rect 247 -2719 261 -2685
rect 189 -2739 261 -2719
rect 535 -2685 607 -2519
rect 535 -2719 549 -2685
rect 583 -2719 607 -2685
rect 535 -2739 607 -2719
rect 189 -2753 607 -2739
rect 189 -2787 213 -2753
rect 247 -2787 281 -2753
rect 315 -2787 481 -2753
rect 515 -2787 549 -2753
rect 583 -2787 607 -2753
rect 189 -2811 607 -2787
rect 1189 -2417 1607 -2393
rect 1189 -2451 1213 -2417
rect 1247 -2451 1281 -2417
rect 1315 -2451 1481 -2417
rect 1515 -2451 1549 -2417
rect 1583 -2451 1607 -2417
rect 1189 -2465 1607 -2451
rect 1189 -2485 1261 -2465
rect 1189 -2519 1213 -2485
rect 1247 -2519 1261 -2485
rect 1189 -2685 1261 -2519
rect 1535 -2485 1607 -2465
rect 1535 -2519 1549 -2485
rect 1583 -2519 1607 -2485
rect 1189 -2719 1213 -2685
rect 1247 -2719 1261 -2685
rect 1189 -2739 1261 -2719
rect 1535 -2685 1607 -2519
rect 1535 -2719 1549 -2685
rect 1583 -2719 1607 -2685
rect 1535 -2739 1607 -2719
rect 1189 -2753 1607 -2739
rect 1189 -2787 1213 -2753
rect 1247 -2787 1281 -2753
rect 1315 -2787 1481 -2753
rect 1515 -2787 1549 -2753
rect 1583 -2787 1607 -2753
rect 1189 -2811 1607 -2787
<< psubdiffcont >>
rect -3940 1702 -3906 1736
rect -3872 1702 -3838 1736
rect -3804 1702 -3770 1736
rect -3736 1702 -3702 1736
rect -3502 1702 -3468 1736
rect -3434 1702 -3400 1736
rect -3366 1702 -3332 1736
rect -3298 1702 -3264 1736
rect -3940 1634 -3906 1668
rect -3298 1634 -3264 1668
rect -3940 1566 -3906 1600
rect -3940 1498 -3906 1532
rect -3940 1264 -3906 1298
rect -3940 1196 -3906 1230
rect -3298 1566 -3264 1600
rect -3298 1498 -3264 1532
rect -3298 1264 -3264 1298
rect -3298 1196 -3264 1230
rect -3940 1128 -3906 1162
rect -3298 1128 -3264 1162
rect -3940 1060 -3906 1094
rect -3872 1060 -3838 1094
rect -3804 1060 -3770 1094
rect -3736 1060 -3702 1094
rect -3502 1060 -3468 1094
rect -3434 1060 -3400 1094
rect -3366 1060 -3332 1094
rect -3298 1060 -3264 1094
rect -2940 1702 -2906 1736
rect -2872 1702 -2838 1736
rect -2804 1702 -2770 1736
rect -2736 1702 -2702 1736
rect -2502 1702 -2468 1736
rect -2434 1702 -2400 1736
rect -2366 1702 -2332 1736
rect -2298 1702 -2264 1736
rect -2940 1634 -2906 1668
rect -2298 1634 -2264 1668
rect -2940 1566 -2906 1600
rect -2940 1498 -2906 1532
rect -2940 1264 -2906 1298
rect -2940 1196 -2906 1230
rect -2298 1566 -2264 1600
rect -2298 1498 -2264 1532
rect -2298 1264 -2264 1298
rect -2298 1196 -2264 1230
rect -2940 1128 -2906 1162
rect -2298 1128 -2264 1162
rect -2940 1060 -2906 1094
rect -2872 1060 -2838 1094
rect -2804 1060 -2770 1094
rect -2736 1060 -2702 1094
rect -2502 1060 -2468 1094
rect -2434 1060 -2400 1094
rect -2366 1060 -2332 1094
rect -2298 1060 -2264 1094
rect -1940 1702 -1906 1736
rect -1872 1702 -1838 1736
rect -1804 1702 -1770 1736
rect -1736 1702 -1702 1736
rect -1502 1702 -1468 1736
rect -1434 1702 -1400 1736
rect -1366 1702 -1332 1736
rect -1298 1702 -1264 1736
rect -1940 1634 -1906 1668
rect -1298 1634 -1264 1668
rect -1940 1566 -1906 1600
rect -1940 1498 -1906 1532
rect -1940 1264 -1906 1298
rect -1940 1196 -1906 1230
rect -1298 1566 -1264 1600
rect -1298 1498 -1264 1532
rect -1298 1264 -1264 1298
rect -1298 1196 -1264 1230
rect -1940 1128 -1906 1162
rect -1298 1128 -1264 1162
rect -1940 1060 -1906 1094
rect -1872 1060 -1838 1094
rect -1804 1060 -1770 1094
rect -1736 1060 -1702 1094
rect -1502 1060 -1468 1094
rect -1434 1060 -1400 1094
rect -1366 1060 -1332 1094
rect -1298 1060 -1264 1094
rect -940 1702 -906 1736
rect -872 1702 -838 1736
rect -804 1702 -770 1736
rect -736 1702 -702 1736
rect -502 1702 -468 1736
rect -434 1702 -400 1736
rect -366 1702 -332 1736
rect -298 1702 -264 1736
rect -940 1634 -906 1668
rect -298 1634 -264 1668
rect -940 1566 -906 1600
rect -940 1498 -906 1532
rect -940 1264 -906 1298
rect -940 1196 -906 1230
rect -298 1566 -264 1600
rect -298 1498 -264 1532
rect -298 1264 -264 1298
rect -298 1196 -264 1230
rect -940 1128 -906 1162
rect -298 1128 -264 1162
rect -940 1060 -906 1094
rect -872 1060 -838 1094
rect -804 1060 -770 1094
rect -736 1060 -702 1094
rect -502 1060 -468 1094
rect -434 1060 -400 1094
rect -366 1060 -332 1094
rect -298 1060 -264 1094
rect 60 1702 94 1736
rect 128 1702 162 1736
rect 196 1702 230 1736
rect 264 1702 298 1736
rect 498 1702 532 1736
rect 566 1702 600 1736
rect 634 1702 668 1736
rect 702 1702 736 1736
rect 60 1634 94 1668
rect 702 1634 736 1668
rect 60 1566 94 1600
rect 60 1498 94 1532
rect 60 1264 94 1298
rect 60 1196 94 1230
rect 702 1566 736 1600
rect 702 1498 736 1532
rect 702 1264 736 1298
rect 702 1196 736 1230
rect 60 1128 94 1162
rect 702 1128 736 1162
rect 60 1060 94 1094
rect 128 1060 162 1094
rect 196 1060 230 1094
rect 264 1060 298 1094
rect 498 1060 532 1094
rect 566 1060 600 1094
rect 634 1060 668 1094
rect 702 1060 736 1094
rect 1060 1702 1094 1736
rect 1128 1702 1162 1736
rect 1196 1702 1230 1736
rect 1264 1702 1298 1736
rect 1498 1702 1532 1736
rect 1566 1702 1600 1736
rect 1634 1702 1668 1736
rect 1702 1702 1736 1736
rect 1060 1634 1094 1668
rect 1702 1634 1736 1668
rect 1060 1566 1094 1600
rect 1060 1498 1094 1532
rect 1060 1264 1094 1298
rect 1060 1196 1094 1230
rect 1702 1566 1736 1600
rect 1702 1498 1736 1532
rect 1702 1264 1736 1298
rect 1702 1196 1736 1230
rect 1060 1128 1094 1162
rect 1702 1128 1736 1162
rect 1060 1060 1094 1094
rect 1128 1060 1162 1094
rect 1196 1060 1230 1094
rect 1264 1060 1298 1094
rect 1498 1060 1532 1094
rect 1566 1060 1600 1094
rect 1634 1060 1668 1094
rect 1702 1060 1736 1094
rect -3940 702 -3906 736
rect -3872 702 -3838 736
rect -3804 702 -3770 736
rect -3736 702 -3702 736
rect -3502 702 -3468 736
rect -3434 702 -3400 736
rect -3366 702 -3332 736
rect -3298 702 -3264 736
rect -3940 634 -3906 668
rect -3298 634 -3264 668
rect -3940 566 -3906 600
rect -3940 498 -3906 532
rect -3940 264 -3906 298
rect -3940 196 -3906 230
rect -3298 566 -3264 600
rect -3298 498 -3264 532
rect -3298 264 -3264 298
rect -3298 196 -3264 230
rect -3940 128 -3906 162
rect -3298 128 -3264 162
rect -3940 60 -3906 94
rect -3872 60 -3838 94
rect -3804 60 -3770 94
rect -3736 60 -3702 94
rect -3502 60 -3468 94
rect -3434 60 -3400 94
rect -3366 60 -3332 94
rect -3298 60 -3264 94
rect -2940 702 -2906 736
rect -2872 702 -2838 736
rect -2804 702 -2770 736
rect -2736 702 -2702 736
rect -2502 702 -2468 736
rect -2434 702 -2400 736
rect -2366 702 -2332 736
rect -2298 702 -2264 736
rect -2940 634 -2906 668
rect -2298 634 -2264 668
rect -2940 566 -2906 600
rect -2940 498 -2906 532
rect -2940 264 -2906 298
rect -2940 196 -2906 230
rect -2298 566 -2264 600
rect -2298 498 -2264 532
rect -2298 264 -2264 298
rect -2298 196 -2264 230
rect -2940 128 -2906 162
rect -2298 128 -2264 162
rect -2940 60 -2906 94
rect -2872 60 -2838 94
rect -2804 60 -2770 94
rect -2736 60 -2702 94
rect -2502 60 -2468 94
rect -2434 60 -2400 94
rect -2366 60 -2332 94
rect -2298 60 -2264 94
rect -1940 702 -1906 736
rect -1872 702 -1838 736
rect -1804 702 -1770 736
rect -1736 702 -1702 736
rect -1502 702 -1468 736
rect -1434 702 -1400 736
rect -1366 702 -1332 736
rect -1298 702 -1264 736
rect -1940 634 -1906 668
rect -1298 634 -1264 668
rect -1940 566 -1906 600
rect -1940 498 -1906 532
rect -1940 264 -1906 298
rect -1940 196 -1906 230
rect -1298 566 -1264 600
rect -1298 498 -1264 532
rect -1298 264 -1264 298
rect -1298 196 -1264 230
rect -1940 128 -1906 162
rect -1298 128 -1264 162
rect -1940 60 -1906 94
rect -1872 60 -1838 94
rect -1804 60 -1770 94
rect -1736 60 -1702 94
rect -1502 60 -1468 94
rect -1434 60 -1400 94
rect -1366 60 -1332 94
rect -1298 60 -1264 94
rect -940 702 -906 736
rect -872 702 -838 736
rect -804 702 -770 736
rect -736 702 -702 736
rect -502 702 -468 736
rect -434 702 -400 736
rect -366 702 -332 736
rect -298 702 -264 736
rect -940 634 -906 668
rect -298 634 -264 668
rect -940 566 -906 600
rect -940 498 -906 532
rect -940 264 -906 298
rect -940 196 -906 230
rect -298 566 -264 600
rect -298 498 -264 532
rect -298 264 -264 298
rect -298 196 -264 230
rect -940 128 -906 162
rect -298 128 -264 162
rect -940 60 -906 94
rect -872 60 -838 94
rect -804 60 -770 94
rect -736 60 -702 94
rect -502 60 -468 94
rect -434 60 -400 94
rect -366 60 -332 94
rect -298 60 -264 94
rect 60 702 94 736
rect 128 702 162 736
rect 196 702 230 736
rect 264 702 298 736
rect 498 702 532 736
rect 566 702 600 736
rect 634 702 668 736
rect 702 702 736 736
rect 60 634 94 668
rect 702 634 736 668
rect 60 566 94 600
rect 60 498 94 532
rect 60 264 94 298
rect 60 196 94 230
rect 702 566 736 600
rect 702 498 736 532
rect 702 264 736 298
rect 702 196 736 230
rect 60 128 94 162
rect 702 128 736 162
rect 60 60 94 94
rect 128 60 162 94
rect 196 60 230 94
rect 264 60 298 94
rect 498 60 532 94
rect 566 60 600 94
rect 634 60 668 94
rect 702 60 736 94
rect 1060 702 1094 736
rect 1128 702 1162 736
rect 1196 702 1230 736
rect 1264 702 1298 736
rect 1498 702 1532 736
rect 1566 702 1600 736
rect 1634 702 1668 736
rect 1702 702 1736 736
rect 1060 634 1094 668
rect 1702 634 1736 668
rect 1060 566 1094 600
rect 1060 498 1094 532
rect 1060 264 1094 298
rect 1060 196 1094 230
rect 1702 566 1736 600
rect 1702 498 1736 532
rect 1702 264 1736 298
rect 1702 196 1736 230
rect 1060 128 1094 162
rect 1702 128 1736 162
rect 1060 60 1094 94
rect 1128 60 1162 94
rect 1196 60 1230 94
rect 1264 60 1298 94
rect 1498 60 1532 94
rect 1566 60 1600 94
rect 1634 60 1668 94
rect 1702 60 1736 94
rect -3940 -298 -3906 -264
rect -3872 -298 -3838 -264
rect -3804 -298 -3770 -264
rect -3736 -298 -3702 -264
rect -3502 -298 -3468 -264
rect -3434 -298 -3400 -264
rect -3366 -298 -3332 -264
rect -3298 -298 -3264 -264
rect -3940 -366 -3906 -332
rect -3298 -366 -3264 -332
rect -3940 -434 -3906 -400
rect -3940 -502 -3906 -468
rect -3940 -736 -3906 -702
rect -3940 -804 -3906 -770
rect -3298 -434 -3264 -400
rect -3298 -502 -3264 -468
rect -3298 -736 -3264 -702
rect -3298 -804 -3264 -770
rect -3940 -872 -3906 -838
rect -3298 -872 -3264 -838
rect -3940 -940 -3906 -906
rect -3872 -940 -3838 -906
rect -3804 -940 -3770 -906
rect -3736 -940 -3702 -906
rect -3502 -940 -3468 -906
rect -3434 -940 -3400 -906
rect -3366 -940 -3332 -906
rect -3298 -940 -3264 -906
rect -2940 -298 -2906 -264
rect -2872 -298 -2838 -264
rect -2804 -298 -2770 -264
rect -2736 -298 -2702 -264
rect -2502 -298 -2468 -264
rect -2434 -298 -2400 -264
rect -2366 -298 -2332 -264
rect -2298 -298 -2264 -264
rect -2940 -366 -2906 -332
rect -2298 -366 -2264 -332
rect -2940 -434 -2906 -400
rect -2940 -502 -2906 -468
rect -2940 -736 -2906 -702
rect -2940 -804 -2906 -770
rect -2298 -434 -2264 -400
rect -2298 -502 -2264 -468
rect -2298 -736 -2264 -702
rect -2298 -804 -2264 -770
rect -2940 -872 -2906 -838
rect -2298 -872 -2264 -838
rect -2940 -940 -2906 -906
rect -2872 -940 -2838 -906
rect -2804 -940 -2770 -906
rect -2736 -940 -2702 -906
rect -2502 -940 -2468 -906
rect -2434 -940 -2400 -906
rect -2366 -940 -2332 -906
rect -2298 -940 -2264 -906
rect -1940 -298 -1906 -264
rect -1872 -298 -1838 -264
rect -1804 -298 -1770 -264
rect -1736 -298 -1702 -264
rect -1502 -298 -1468 -264
rect -1434 -298 -1400 -264
rect -1366 -298 -1332 -264
rect -1298 -298 -1264 -264
rect -1940 -366 -1906 -332
rect -1298 -366 -1264 -332
rect -1940 -434 -1906 -400
rect -1940 -502 -1906 -468
rect -1940 -736 -1906 -702
rect -1940 -804 -1906 -770
rect -1298 -434 -1264 -400
rect -1298 -502 -1264 -468
rect -1298 -736 -1264 -702
rect -1298 -804 -1264 -770
rect -1940 -872 -1906 -838
rect -1298 -872 -1264 -838
rect -1940 -940 -1906 -906
rect -1872 -940 -1838 -906
rect -1804 -940 -1770 -906
rect -1736 -940 -1702 -906
rect -1502 -940 -1468 -906
rect -1434 -940 -1400 -906
rect -1366 -940 -1332 -906
rect -1298 -940 -1264 -906
rect -940 -298 -906 -264
rect -872 -298 -838 -264
rect -804 -298 -770 -264
rect -736 -298 -702 -264
rect -502 -298 -468 -264
rect -434 -298 -400 -264
rect -366 -298 -332 -264
rect -298 -298 -264 -264
rect -940 -366 -906 -332
rect -298 -366 -264 -332
rect -940 -434 -906 -400
rect -940 -502 -906 -468
rect -940 -736 -906 -702
rect -940 -804 -906 -770
rect -298 -434 -264 -400
rect -298 -502 -264 -468
rect -298 -736 -264 -702
rect -298 -804 -264 -770
rect -940 -872 -906 -838
rect -298 -872 -264 -838
rect -940 -940 -906 -906
rect -872 -940 -838 -906
rect -804 -940 -770 -906
rect -736 -940 -702 -906
rect -502 -940 -468 -906
rect -434 -940 -400 -906
rect -366 -940 -332 -906
rect -298 -940 -264 -906
rect 60 -298 94 -264
rect 128 -298 162 -264
rect 196 -298 230 -264
rect 264 -298 298 -264
rect 498 -298 532 -264
rect 566 -298 600 -264
rect 634 -298 668 -264
rect 702 -298 736 -264
rect 60 -366 94 -332
rect 702 -366 736 -332
rect 60 -434 94 -400
rect 60 -502 94 -468
rect 60 -736 94 -702
rect 60 -804 94 -770
rect 702 -434 736 -400
rect 702 -502 736 -468
rect 702 -736 736 -702
rect 702 -804 736 -770
rect 60 -872 94 -838
rect 702 -872 736 -838
rect 60 -940 94 -906
rect 128 -940 162 -906
rect 196 -940 230 -906
rect 264 -940 298 -906
rect 498 -940 532 -906
rect 566 -940 600 -906
rect 634 -940 668 -906
rect 702 -940 736 -906
rect 1060 -298 1094 -264
rect 1128 -298 1162 -264
rect 1196 -298 1230 -264
rect 1264 -298 1298 -264
rect 1498 -298 1532 -264
rect 1566 -298 1600 -264
rect 1634 -298 1668 -264
rect 1702 -298 1736 -264
rect 1060 -366 1094 -332
rect 1702 -366 1736 -332
rect 1060 -434 1094 -400
rect 1060 -502 1094 -468
rect 1060 -736 1094 -702
rect 1060 -804 1094 -770
rect 1702 -434 1736 -400
rect 1702 -502 1736 -468
rect 1702 -736 1736 -702
rect 1702 -804 1736 -770
rect 1060 -872 1094 -838
rect 1702 -872 1736 -838
rect 1060 -940 1094 -906
rect 1128 -940 1162 -906
rect 1196 -940 1230 -906
rect 1264 -940 1298 -906
rect 1498 -940 1532 -906
rect 1566 -940 1600 -906
rect 1634 -940 1668 -906
rect 1702 -940 1736 -906
rect -3940 -1298 -3906 -1264
rect -3872 -1298 -3838 -1264
rect -3804 -1298 -3770 -1264
rect -3736 -1298 -3702 -1264
rect -3502 -1298 -3468 -1264
rect -3434 -1298 -3400 -1264
rect -3366 -1298 -3332 -1264
rect -3298 -1298 -3264 -1264
rect -3940 -1366 -3906 -1332
rect -3298 -1366 -3264 -1332
rect -3940 -1434 -3906 -1400
rect -3940 -1502 -3906 -1468
rect -3940 -1736 -3906 -1702
rect -3940 -1804 -3906 -1770
rect -3298 -1434 -3264 -1400
rect -3298 -1502 -3264 -1468
rect -3298 -1736 -3264 -1702
rect -3298 -1804 -3264 -1770
rect -3940 -1872 -3906 -1838
rect -3298 -1872 -3264 -1838
rect -3940 -1940 -3906 -1906
rect -3872 -1940 -3838 -1906
rect -3804 -1940 -3770 -1906
rect -3736 -1940 -3702 -1906
rect -3502 -1940 -3468 -1906
rect -3434 -1940 -3400 -1906
rect -3366 -1940 -3332 -1906
rect -3298 -1940 -3264 -1906
rect -2940 -1298 -2906 -1264
rect -2872 -1298 -2838 -1264
rect -2804 -1298 -2770 -1264
rect -2736 -1298 -2702 -1264
rect -2502 -1298 -2468 -1264
rect -2434 -1298 -2400 -1264
rect -2366 -1298 -2332 -1264
rect -2298 -1298 -2264 -1264
rect -2940 -1366 -2906 -1332
rect -2298 -1366 -2264 -1332
rect -2940 -1434 -2906 -1400
rect -2940 -1502 -2906 -1468
rect -2940 -1736 -2906 -1702
rect -2940 -1804 -2906 -1770
rect -2298 -1434 -2264 -1400
rect -2298 -1502 -2264 -1468
rect -2298 -1736 -2264 -1702
rect -2298 -1804 -2264 -1770
rect -2940 -1872 -2906 -1838
rect -2298 -1872 -2264 -1838
rect -2940 -1940 -2906 -1906
rect -2872 -1940 -2838 -1906
rect -2804 -1940 -2770 -1906
rect -2736 -1940 -2702 -1906
rect -2502 -1940 -2468 -1906
rect -2434 -1940 -2400 -1906
rect -2366 -1940 -2332 -1906
rect -2298 -1940 -2264 -1906
rect -1940 -1298 -1906 -1264
rect -1872 -1298 -1838 -1264
rect -1804 -1298 -1770 -1264
rect -1736 -1298 -1702 -1264
rect -1502 -1298 -1468 -1264
rect -1434 -1298 -1400 -1264
rect -1366 -1298 -1332 -1264
rect -1298 -1298 -1264 -1264
rect -1940 -1366 -1906 -1332
rect -1298 -1366 -1264 -1332
rect -1940 -1434 -1906 -1400
rect -1940 -1502 -1906 -1468
rect -1940 -1736 -1906 -1702
rect -1940 -1804 -1906 -1770
rect -1298 -1434 -1264 -1400
rect -1298 -1502 -1264 -1468
rect -1298 -1736 -1264 -1702
rect -1298 -1804 -1264 -1770
rect -1940 -1872 -1906 -1838
rect -1298 -1872 -1264 -1838
rect -1940 -1940 -1906 -1906
rect -1872 -1940 -1838 -1906
rect -1804 -1940 -1770 -1906
rect -1736 -1940 -1702 -1906
rect -1502 -1940 -1468 -1906
rect -1434 -1940 -1400 -1906
rect -1366 -1940 -1332 -1906
rect -1298 -1940 -1264 -1906
rect -940 -1298 -906 -1264
rect -872 -1298 -838 -1264
rect -804 -1298 -770 -1264
rect -736 -1298 -702 -1264
rect -502 -1298 -468 -1264
rect -434 -1298 -400 -1264
rect -366 -1298 -332 -1264
rect -298 -1298 -264 -1264
rect -940 -1366 -906 -1332
rect -298 -1366 -264 -1332
rect -940 -1434 -906 -1400
rect -940 -1502 -906 -1468
rect -940 -1736 -906 -1702
rect -940 -1804 -906 -1770
rect -298 -1434 -264 -1400
rect -298 -1502 -264 -1468
rect -298 -1736 -264 -1702
rect -298 -1804 -264 -1770
rect -940 -1872 -906 -1838
rect -298 -1872 -264 -1838
rect -940 -1940 -906 -1906
rect -872 -1940 -838 -1906
rect -804 -1940 -770 -1906
rect -736 -1940 -702 -1906
rect -502 -1940 -468 -1906
rect -434 -1940 -400 -1906
rect -366 -1940 -332 -1906
rect -298 -1940 -264 -1906
rect 60 -1298 94 -1264
rect 128 -1298 162 -1264
rect 196 -1298 230 -1264
rect 264 -1298 298 -1264
rect 498 -1298 532 -1264
rect 566 -1298 600 -1264
rect 634 -1298 668 -1264
rect 702 -1298 736 -1264
rect 60 -1366 94 -1332
rect 702 -1366 736 -1332
rect 60 -1434 94 -1400
rect 60 -1502 94 -1468
rect 60 -1736 94 -1702
rect 60 -1804 94 -1770
rect 702 -1434 736 -1400
rect 702 -1502 736 -1468
rect 702 -1736 736 -1702
rect 702 -1804 736 -1770
rect 60 -1872 94 -1838
rect 702 -1872 736 -1838
rect 60 -1940 94 -1906
rect 128 -1940 162 -1906
rect 196 -1940 230 -1906
rect 264 -1940 298 -1906
rect 498 -1940 532 -1906
rect 566 -1940 600 -1906
rect 634 -1940 668 -1906
rect 702 -1940 736 -1906
rect 1060 -1298 1094 -1264
rect 1128 -1298 1162 -1264
rect 1196 -1298 1230 -1264
rect 1264 -1298 1298 -1264
rect 1498 -1298 1532 -1264
rect 1566 -1298 1600 -1264
rect 1634 -1298 1668 -1264
rect 1702 -1298 1736 -1264
rect 1060 -1366 1094 -1332
rect 1702 -1366 1736 -1332
rect 1060 -1434 1094 -1400
rect 1060 -1502 1094 -1468
rect 1060 -1736 1094 -1702
rect 1060 -1804 1094 -1770
rect 1702 -1434 1736 -1400
rect 1702 -1502 1736 -1468
rect 1702 -1736 1736 -1702
rect 1702 -1804 1736 -1770
rect 1060 -1872 1094 -1838
rect 1702 -1872 1736 -1838
rect 1060 -1940 1094 -1906
rect 1128 -1940 1162 -1906
rect 1196 -1940 1230 -1906
rect 1264 -1940 1298 -1906
rect 1498 -1940 1532 -1906
rect 1566 -1940 1600 -1906
rect 1634 -1940 1668 -1906
rect 1702 -1940 1736 -1906
rect -3940 -2298 -3906 -2264
rect -3872 -2298 -3838 -2264
rect -3804 -2298 -3770 -2264
rect -3736 -2298 -3702 -2264
rect -3502 -2298 -3468 -2264
rect -3434 -2298 -3400 -2264
rect -3366 -2298 -3332 -2264
rect -3298 -2298 -3264 -2264
rect -3940 -2366 -3906 -2332
rect -3298 -2366 -3264 -2332
rect -3940 -2434 -3906 -2400
rect -3940 -2502 -3906 -2468
rect -3940 -2736 -3906 -2702
rect -3940 -2804 -3906 -2770
rect -3298 -2434 -3264 -2400
rect -3298 -2502 -3264 -2468
rect -3298 -2736 -3264 -2702
rect -3298 -2804 -3264 -2770
rect -3940 -2872 -3906 -2838
rect -3298 -2872 -3264 -2838
rect -3940 -2940 -3906 -2906
rect -3872 -2940 -3838 -2906
rect -3804 -2940 -3770 -2906
rect -3736 -2940 -3702 -2906
rect -3502 -2940 -3468 -2906
rect -3434 -2940 -3400 -2906
rect -3366 -2940 -3332 -2906
rect -3298 -2940 -3264 -2906
rect -2940 -2298 -2906 -2264
rect -2872 -2298 -2838 -2264
rect -2804 -2298 -2770 -2264
rect -2736 -2298 -2702 -2264
rect -2502 -2298 -2468 -2264
rect -2434 -2298 -2400 -2264
rect -2366 -2298 -2332 -2264
rect -2298 -2298 -2264 -2264
rect -2940 -2366 -2906 -2332
rect -2298 -2366 -2264 -2332
rect -2940 -2434 -2906 -2400
rect -2940 -2502 -2906 -2468
rect -2940 -2736 -2906 -2702
rect -2940 -2804 -2906 -2770
rect -2298 -2434 -2264 -2400
rect -2298 -2502 -2264 -2468
rect -2298 -2736 -2264 -2702
rect -2298 -2804 -2264 -2770
rect -2940 -2872 -2906 -2838
rect -2298 -2872 -2264 -2838
rect -2940 -2940 -2906 -2906
rect -2872 -2940 -2838 -2906
rect -2804 -2940 -2770 -2906
rect -2736 -2940 -2702 -2906
rect -2502 -2940 -2468 -2906
rect -2434 -2940 -2400 -2906
rect -2366 -2940 -2332 -2906
rect -2298 -2940 -2264 -2906
rect -1940 -2298 -1906 -2264
rect -1872 -2298 -1838 -2264
rect -1804 -2298 -1770 -2264
rect -1736 -2298 -1702 -2264
rect -1502 -2298 -1468 -2264
rect -1434 -2298 -1400 -2264
rect -1366 -2298 -1332 -2264
rect -1298 -2298 -1264 -2264
rect -1940 -2366 -1906 -2332
rect -1298 -2366 -1264 -2332
rect -1940 -2434 -1906 -2400
rect -1940 -2502 -1906 -2468
rect -1940 -2736 -1906 -2702
rect -1940 -2804 -1906 -2770
rect -1298 -2434 -1264 -2400
rect -1298 -2502 -1264 -2468
rect -1298 -2736 -1264 -2702
rect -1298 -2804 -1264 -2770
rect -1940 -2872 -1906 -2838
rect -1298 -2872 -1264 -2838
rect -1940 -2940 -1906 -2906
rect -1872 -2940 -1838 -2906
rect -1804 -2940 -1770 -2906
rect -1736 -2940 -1702 -2906
rect -1502 -2940 -1468 -2906
rect -1434 -2940 -1400 -2906
rect -1366 -2940 -1332 -2906
rect -1298 -2940 -1264 -2906
rect -940 -2298 -906 -2264
rect -872 -2298 -838 -2264
rect -804 -2298 -770 -2264
rect -736 -2298 -702 -2264
rect -502 -2298 -468 -2264
rect -434 -2298 -400 -2264
rect -366 -2298 -332 -2264
rect -298 -2298 -264 -2264
rect -940 -2366 -906 -2332
rect -298 -2366 -264 -2332
rect -940 -2434 -906 -2400
rect -940 -2502 -906 -2468
rect -940 -2736 -906 -2702
rect -940 -2804 -906 -2770
rect -298 -2434 -264 -2400
rect -298 -2502 -264 -2468
rect -298 -2736 -264 -2702
rect -298 -2804 -264 -2770
rect -940 -2872 -906 -2838
rect -298 -2872 -264 -2838
rect -940 -2940 -906 -2906
rect -872 -2940 -838 -2906
rect -804 -2940 -770 -2906
rect -736 -2940 -702 -2906
rect -502 -2940 -468 -2906
rect -434 -2940 -400 -2906
rect -366 -2940 -332 -2906
rect -298 -2940 -264 -2906
rect 60 -2298 94 -2264
rect 128 -2298 162 -2264
rect 196 -2298 230 -2264
rect 264 -2298 298 -2264
rect 498 -2298 532 -2264
rect 566 -2298 600 -2264
rect 634 -2298 668 -2264
rect 702 -2298 736 -2264
rect 60 -2366 94 -2332
rect 702 -2366 736 -2332
rect 60 -2434 94 -2400
rect 60 -2502 94 -2468
rect 60 -2736 94 -2702
rect 60 -2804 94 -2770
rect 702 -2434 736 -2400
rect 702 -2502 736 -2468
rect 702 -2736 736 -2702
rect 702 -2804 736 -2770
rect 60 -2872 94 -2838
rect 702 -2872 736 -2838
rect 60 -2940 94 -2906
rect 128 -2940 162 -2906
rect 196 -2940 230 -2906
rect 264 -2940 298 -2906
rect 498 -2940 532 -2906
rect 566 -2940 600 -2906
rect 634 -2940 668 -2906
rect 702 -2940 736 -2906
rect 1060 -2298 1094 -2264
rect 1128 -2298 1162 -2264
rect 1196 -2298 1230 -2264
rect 1264 -2298 1298 -2264
rect 1498 -2298 1532 -2264
rect 1566 -2298 1600 -2264
rect 1634 -2298 1668 -2264
rect 1702 -2298 1736 -2264
rect 1060 -2366 1094 -2332
rect 1702 -2366 1736 -2332
rect 1060 -2434 1094 -2400
rect 1060 -2502 1094 -2468
rect 1060 -2736 1094 -2702
rect 1060 -2804 1094 -2770
rect 1702 -2434 1736 -2400
rect 1702 -2502 1736 -2468
rect 1702 -2736 1736 -2702
rect 1702 -2804 1736 -2770
rect 1060 -2872 1094 -2838
rect 1702 -2872 1736 -2838
rect 1060 -2940 1094 -2906
rect 1128 -2940 1162 -2906
rect 1196 -2940 1230 -2906
rect 1264 -2940 1298 -2906
rect 1498 -2940 1532 -2906
rect 1566 -2940 1600 -2906
rect 1634 -2940 1668 -2906
rect 1702 -2940 1736 -2906
<< nsubdiffcont >>
rect -3787 1549 -3753 1583
rect -3719 1549 -3685 1583
rect -3519 1549 -3485 1583
rect -3451 1549 -3417 1583
rect -3787 1481 -3753 1515
rect -3451 1481 -3417 1515
rect -3787 1281 -3753 1315
rect -3451 1281 -3417 1315
rect -3787 1213 -3753 1247
rect -3719 1213 -3685 1247
rect -3519 1213 -3485 1247
rect -3451 1213 -3417 1247
rect -2787 1549 -2753 1583
rect -2719 1549 -2685 1583
rect -2519 1549 -2485 1583
rect -2451 1549 -2417 1583
rect -2787 1481 -2753 1515
rect -2451 1481 -2417 1515
rect -2787 1281 -2753 1315
rect -2451 1281 -2417 1315
rect -2787 1213 -2753 1247
rect -2719 1213 -2685 1247
rect -2519 1213 -2485 1247
rect -2451 1213 -2417 1247
rect -1787 1549 -1753 1583
rect -1719 1549 -1685 1583
rect -1519 1549 -1485 1583
rect -1451 1549 -1417 1583
rect -1787 1481 -1753 1515
rect -1451 1481 -1417 1515
rect -1787 1281 -1753 1315
rect -1451 1281 -1417 1315
rect -1787 1213 -1753 1247
rect -1719 1213 -1685 1247
rect -1519 1213 -1485 1247
rect -1451 1213 -1417 1247
rect -787 1549 -753 1583
rect -719 1549 -685 1583
rect -519 1549 -485 1583
rect -451 1549 -417 1583
rect -787 1481 -753 1515
rect -451 1481 -417 1515
rect -787 1281 -753 1315
rect -451 1281 -417 1315
rect -787 1213 -753 1247
rect -719 1213 -685 1247
rect -519 1213 -485 1247
rect -451 1213 -417 1247
rect 213 1549 247 1583
rect 281 1549 315 1583
rect 481 1549 515 1583
rect 549 1549 583 1583
rect 213 1481 247 1515
rect 549 1481 583 1515
rect 213 1281 247 1315
rect 549 1281 583 1315
rect 213 1213 247 1247
rect 281 1213 315 1247
rect 481 1213 515 1247
rect 549 1213 583 1247
rect 1213 1549 1247 1583
rect 1281 1549 1315 1583
rect 1481 1549 1515 1583
rect 1549 1549 1583 1583
rect 1213 1481 1247 1515
rect 1549 1481 1583 1515
rect 1213 1281 1247 1315
rect 1549 1281 1583 1315
rect 1213 1213 1247 1247
rect 1281 1213 1315 1247
rect 1481 1213 1515 1247
rect 1549 1213 1583 1247
rect -3787 549 -3753 583
rect -3719 549 -3685 583
rect -3519 549 -3485 583
rect -3451 549 -3417 583
rect -3787 481 -3753 515
rect -3451 481 -3417 515
rect -3787 281 -3753 315
rect -3451 281 -3417 315
rect -3787 213 -3753 247
rect -3719 213 -3685 247
rect -3519 213 -3485 247
rect -3451 213 -3417 247
rect -2787 549 -2753 583
rect -2719 549 -2685 583
rect -2519 549 -2485 583
rect -2451 549 -2417 583
rect -2787 481 -2753 515
rect -2451 481 -2417 515
rect -2787 281 -2753 315
rect -2451 281 -2417 315
rect -2787 213 -2753 247
rect -2719 213 -2685 247
rect -2519 213 -2485 247
rect -2451 213 -2417 247
rect -1787 549 -1753 583
rect -1719 549 -1685 583
rect -1519 549 -1485 583
rect -1451 549 -1417 583
rect -1787 481 -1753 515
rect -1451 481 -1417 515
rect -1787 281 -1753 315
rect -1451 281 -1417 315
rect -1787 213 -1753 247
rect -1719 213 -1685 247
rect -1519 213 -1485 247
rect -1451 213 -1417 247
rect -787 549 -753 583
rect -719 549 -685 583
rect -519 549 -485 583
rect -451 549 -417 583
rect -787 481 -753 515
rect -451 481 -417 515
rect -787 281 -753 315
rect -451 281 -417 315
rect -787 213 -753 247
rect -719 213 -685 247
rect -519 213 -485 247
rect -451 213 -417 247
rect 213 549 247 583
rect 281 549 315 583
rect 481 549 515 583
rect 549 549 583 583
rect 213 481 247 515
rect 549 481 583 515
rect 213 281 247 315
rect 549 281 583 315
rect 213 213 247 247
rect 281 213 315 247
rect 481 213 515 247
rect 549 213 583 247
rect 1213 549 1247 583
rect 1281 549 1315 583
rect 1481 549 1515 583
rect 1549 549 1583 583
rect 1213 481 1247 515
rect 1549 481 1583 515
rect 1213 281 1247 315
rect 1549 281 1583 315
rect 1213 213 1247 247
rect 1281 213 1315 247
rect 1481 213 1515 247
rect 1549 213 1583 247
rect -3787 -451 -3753 -417
rect -3719 -451 -3685 -417
rect -3519 -451 -3485 -417
rect -3451 -451 -3417 -417
rect -3787 -519 -3753 -485
rect -3451 -519 -3417 -485
rect -3787 -719 -3753 -685
rect -3451 -719 -3417 -685
rect -3787 -787 -3753 -753
rect -3719 -787 -3685 -753
rect -3519 -787 -3485 -753
rect -3451 -787 -3417 -753
rect -2787 -451 -2753 -417
rect -2719 -451 -2685 -417
rect -2519 -451 -2485 -417
rect -2451 -451 -2417 -417
rect -2787 -519 -2753 -485
rect -2451 -519 -2417 -485
rect -2787 -719 -2753 -685
rect -2451 -719 -2417 -685
rect -2787 -787 -2753 -753
rect -2719 -787 -2685 -753
rect -2519 -787 -2485 -753
rect -2451 -787 -2417 -753
rect -1787 -451 -1753 -417
rect -1719 -451 -1685 -417
rect -1519 -451 -1485 -417
rect -1451 -451 -1417 -417
rect -1787 -519 -1753 -485
rect -1451 -519 -1417 -485
rect -1787 -719 -1753 -685
rect -1451 -719 -1417 -685
rect -1787 -787 -1753 -753
rect -1719 -787 -1685 -753
rect -1519 -787 -1485 -753
rect -1451 -787 -1417 -753
rect -787 -451 -753 -417
rect -719 -451 -685 -417
rect -519 -451 -485 -417
rect -451 -451 -417 -417
rect -787 -519 -753 -485
rect -451 -519 -417 -485
rect -787 -719 -753 -685
rect -451 -719 -417 -685
rect -787 -787 -753 -753
rect -719 -787 -685 -753
rect -519 -787 -485 -753
rect -451 -787 -417 -753
rect 213 -451 247 -417
rect 281 -451 315 -417
rect 481 -451 515 -417
rect 549 -451 583 -417
rect 213 -519 247 -485
rect 549 -519 583 -485
rect 213 -719 247 -685
rect 549 -719 583 -685
rect 213 -787 247 -753
rect 281 -787 315 -753
rect 481 -787 515 -753
rect 549 -787 583 -753
rect 1213 -451 1247 -417
rect 1281 -451 1315 -417
rect 1481 -451 1515 -417
rect 1549 -451 1583 -417
rect 1213 -519 1247 -485
rect 1549 -519 1583 -485
rect 1213 -719 1247 -685
rect 1549 -719 1583 -685
rect 1213 -787 1247 -753
rect 1281 -787 1315 -753
rect 1481 -787 1515 -753
rect 1549 -787 1583 -753
rect -3787 -1451 -3753 -1417
rect -3719 -1451 -3685 -1417
rect -3519 -1451 -3485 -1417
rect -3451 -1451 -3417 -1417
rect -3787 -1519 -3753 -1485
rect -3451 -1519 -3417 -1485
rect -3787 -1719 -3753 -1685
rect -3451 -1719 -3417 -1685
rect -3787 -1787 -3753 -1753
rect -3719 -1787 -3685 -1753
rect -3519 -1787 -3485 -1753
rect -3451 -1787 -3417 -1753
rect -2787 -1451 -2753 -1417
rect -2719 -1451 -2685 -1417
rect -2519 -1451 -2485 -1417
rect -2451 -1451 -2417 -1417
rect -2787 -1519 -2753 -1485
rect -2451 -1519 -2417 -1485
rect -2787 -1719 -2753 -1685
rect -2451 -1719 -2417 -1685
rect -2787 -1787 -2753 -1753
rect -2719 -1787 -2685 -1753
rect -2519 -1787 -2485 -1753
rect -2451 -1787 -2417 -1753
rect -1787 -1451 -1753 -1417
rect -1719 -1451 -1685 -1417
rect -1519 -1451 -1485 -1417
rect -1451 -1451 -1417 -1417
rect -1787 -1519 -1753 -1485
rect -1451 -1519 -1417 -1485
rect -1787 -1719 -1753 -1685
rect -1451 -1719 -1417 -1685
rect -1787 -1787 -1753 -1753
rect -1719 -1787 -1685 -1753
rect -1519 -1787 -1485 -1753
rect -1451 -1787 -1417 -1753
rect -787 -1451 -753 -1417
rect -719 -1451 -685 -1417
rect -519 -1451 -485 -1417
rect -451 -1451 -417 -1417
rect -787 -1519 -753 -1485
rect -451 -1519 -417 -1485
rect -787 -1719 -753 -1685
rect -451 -1719 -417 -1685
rect -787 -1787 -753 -1753
rect -719 -1787 -685 -1753
rect -519 -1787 -485 -1753
rect -451 -1787 -417 -1753
rect 213 -1451 247 -1417
rect 281 -1451 315 -1417
rect 481 -1451 515 -1417
rect 549 -1451 583 -1417
rect 213 -1519 247 -1485
rect 549 -1519 583 -1485
rect 213 -1719 247 -1685
rect 549 -1719 583 -1685
rect 213 -1787 247 -1753
rect 281 -1787 315 -1753
rect 481 -1787 515 -1753
rect 549 -1787 583 -1753
rect 1213 -1451 1247 -1417
rect 1281 -1451 1315 -1417
rect 1481 -1451 1515 -1417
rect 1549 -1451 1583 -1417
rect 1213 -1519 1247 -1485
rect 1549 -1519 1583 -1485
rect 1213 -1719 1247 -1685
rect 1549 -1719 1583 -1685
rect 1213 -1787 1247 -1753
rect 1281 -1787 1315 -1753
rect 1481 -1787 1515 -1753
rect 1549 -1787 1583 -1753
rect -3787 -2451 -3753 -2417
rect -3719 -2451 -3685 -2417
rect -3519 -2451 -3485 -2417
rect -3451 -2451 -3417 -2417
rect -3787 -2519 -3753 -2485
rect -3451 -2519 -3417 -2485
rect -3787 -2719 -3753 -2685
rect -3451 -2719 -3417 -2685
rect -3787 -2787 -3753 -2753
rect -3719 -2787 -3685 -2753
rect -3519 -2787 -3485 -2753
rect -3451 -2787 -3417 -2753
rect -2787 -2451 -2753 -2417
rect -2719 -2451 -2685 -2417
rect -2519 -2451 -2485 -2417
rect -2451 -2451 -2417 -2417
rect -2787 -2519 -2753 -2485
rect -2451 -2519 -2417 -2485
rect -2787 -2719 -2753 -2685
rect -2451 -2719 -2417 -2685
rect -2787 -2787 -2753 -2753
rect -2719 -2787 -2685 -2753
rect -2519 -2787 -2485 -2753
rect -2451 -2787 -2417 -2753
rect -1787 -2451 -1753 -2417
rect -1719 -2451 -1685 -2417
rect -1519 -2451 -1485 -2417
rect -1451 -2451 -1417 -2417
rect -1787 -2519 -1753 -2485
rect -1451 -2519 -1417 -2485
rect -1787 -2719 -1753 -2685
rect -1451 -2719 -1417 -2685
rect -1787 -2787 -1753 -2753
rect -1719 -2787 -1685 -2753
rect -1519 -2787 -1485 -2753
rect -1451 -2787 -1417 -2753
rect -787 -2451 -753 -2417
rect -719 -2451 -685 -2417
rect -519 -2451 -485 -2417
rect -451 -2451 -417 -2417
rect -787 -2519 -753 -2485
rect -451 -2519 -417 -2485
rect -787 -2719 -753 -2685
rect -451 -2719 -417 -2685
rect -787 -2787 -753 -2753
rect -719 -2787 -685 -2753
rect -519 -2787 -485 -2753
rect -451 -2787 -417 -2753
rect 213 -2451 247 -2417
rect 281 -2451 315 -2417
rect 481 -2451 515 -2417
rect 549 -2451 583 -2417
rect 213 -2519 247 -2485
rect 549 -2519 583 -2485
rect 213 -2719 247 -2685
rect 549 -2719 583 -2685
rect 213 -2787 247 -2753
rect 281 -2787 315 -2753
rect 481 -2787 515 -2753
rect 549 -2787 583 -2753
rect 1213 -2451 1247 -2417
rect 1281 -2451 1315 -2417
rect 1481 -2451 1515 -2417
rect 1549 -2451 1583 -2417
rect 1213 -2519 1247 -2485
rect 1549 -2519 1583 -2485
rect 1213 -2719 1247 -2685
rect 1549 -2719 1583 -2685
rect 1213 -2787 1247 -2753
rect 1281 -2787 1315 -2753
rect 1481 -2787 1515 -2753
rect 1549 -2787 1583 -2753
<< xpolycontact >>
rect 2250 -2460 2300 -2060
rect -130 -3370 310 -3300
<< locali >>
rect -3974 1736 -3230 1770
rect -3974 1702 -3940 1736
rect -3906 1702 -3872 1736
rect -3838 1702 -3804 1736
rect -3770 1702 -3736 1736
rect -3702 1702 -3502 1736
rect -3468 1702 -3434 1736
rect -3400 1702 -3366 1736
rect -3332 1702 -3298 1736
rect -3264 1702 -3230 1736
rect -3974 1669 -3230 1702
rect -3974 1668 -3873 1669
rect -3974 1634 -3940 1668
rect -3906 1634 -3873 1668
rect -3974 1600 -3873 1634
rect -3331 1668 -3230 1669
rect -3331 1634 -3298 1668
rect -3264 1634 -3230 1668
rect -3974 1566 -3940 1600
rect -3906 1566 -3873 1600
rect -3974 1532 -3873 1566
rect -3974 1498 -3940 1532
rect -3906 1498 -3873 1532
rect -3974 1298 -3873 1498
rect -3974 1264 -3940 1298
rect -3906 1264 -3873 1298
rect -3974 1230 -3873 1264
rect -3974 1196 -3940 1230
rect -3906 1196 -3873 1230
rect -3974 1162 -3873 1196
rect -3811 1583 -3393 1607
rect -3811 1549 -3787 1583
rect -3753 1549 -3719 1583
rect -3685 1549 -3519 1583
rect -3485 1549 -3451 1583
rect -3417 1549 -3393 1583
rect -3811 1535 -3393 1549
rect -3811 1515 -3739 1535
rect -3811 1481 -3787 1515
rect -3753 1481 -3739 1515
rect -3811 1315 -3739 1481
rect -3465 1515 -3393 1535
rect -3465 1481 -3451 1515
rect -3417 1481 -3393 1515
rect -3681 1463 -3523 1477
rect -3681 1429 -3667 1463
rect -3633 1449 -3571 1463
rect -3537 1429 -3523 1463
rect -3681 1367 -3653 1429
rect -3551 1367 -3523 1429
rect -3681 1333 -3667 1367
rect -3633 1333 -3571 1347
rect -3537 1333 -3523 1367
rect -3681 1319 -3523 1333
rect -3811 1281 -3787 1315
rect -3753 1281 -3739 1315
rect -3811 1261 -3739 1281
rect -3465 1315 -3393 1481
rect -3465 1281 -3451 1315
rect -3417 1281 -3393 1315
rect -3465 1261 -3393 1281
rect -3811 1247 -3393 1261
rect -3811 1213 -3787 1247
rect -3753 1213 -3719 1247
rect -3685 1213 -3519 1247
rect -3485 1213 -3451 1247
rect -3417 1213 -3393 1247
rect -3811 1189 -3393 1213
rect -3331 1600 -3230 1634
rect -3331 1566 -3298 1600
rect -3264 1566 -3230 1600
rect -3331 1532 -3230 1566
rect -3331 1498 -3298 1532
rect -3264 1498 -3230 1532
rect -3331 1298 -3230 1498
rect -3331 1264 -3298 1298
rect -3264 1264 -3230 1298
rect -3331 1230 -3230 1264
rect -3331 1196 -3298 1230
rect -3264 1196 -3230 1230
rect -3974 1128 -3940 1162
rect -3906 1128 -3873 1162
rect -3974 1127 -3873 1128
rect -3331 1162 -3230 1196
rect -3331 1128 -3298 1162
rect -3264 1128 -3230 1162
rect -3331 1127 -3230 1128
rect -3974 1094 -3230 1127
rect -3974 1060 -3940 1094
rect -3906 1060 -3872 1094
rect -3838 1060 -3804 1094
rect -3770 1060 -3736 1094
rect -3702 1060 -3502 1094
rect -3468 1060 -3434 1094
rect -3400 1060 -3366 1094
rect -3332 1060 -3298 1094
rect -3264 1060 -3230 1094
rect -3974 1026 -3230 1060
rect -2974 1736 -2230 1770
rect -2974 1702 -2940 1736
rect -2906 1702 -2872 1736
rect -2838 1702 -2804 1736
rect -2770 1702 -2736 1736
rect -2702 1702 -2502 1736
rect -2468 1702 -2434 1736
rect -2400 1702 -2366 1736
rect -2332 1702 -2298 1736
rect -2264 1702 -2230 1736
rect -2974 1669 -2230 1702
rect -2974 1668 -2873 1669
rect -2974 1634 -2940 1668
rect -2906 1634 -2873 1668
rect -2974 1600 -2873 1634
rect -2331 1668 -2230 1669
rect -2331 1634 -2298 1668
rect -2264 1634 -2230 1668
rect -2974 1566 -2940 1600
rect -2906 1566 -2873 1600
rect -2974 1532 -2873 1566
rect -2974 1498 -2940 1532
rect -2906 1498 -2873 1532
rect -2974 1298 -2873 1498
rect -2974 1264 -2940 1298
rect -2906 1264 -2873 1298
rect -2974 1230 -2873 1264
rect -2974 1196 -2940 1230
rect -2906 1196 -2873 1230
rect -2974 1162 -2873 1196
rect -2811 1583 -2393 1607
rect -2811 1549 -2787 1583
rect -2753 1549 -2719 1583
rect -2685 1549 -2519 1583
rect -2485 1549 -2451 1583
rect -2417 1549 -2393 1583
rect -2811 1535 -2393 1549
rect -2811 1515 -2739 1535
rect -2811 1481 -2787 1515
rect -2753 1481 -2739 1515
rect -2811 1315 -2739 1481
rect -2465 1515 -2393 1535
rect -2465 1481 -2451 1515
rect -2417 1481 -2393 1515
rect -2681 1463 -2523 1477
rect -2681 1429 -2667 1463
rect -2633 1449 -2571 1463
rect -2537 1429 -2523 1463
rect -2681 1367 -2653 1429
rect -2551 1367 -2523 1429
rect -2681 1333 -2667 1367
rect -2633 1333 -2571 1347
rect -2537 1333 -2523 1367
rect -2681 1319 -2523 1333
rect -2811 1281 -2787 1315
rect -2753 1281 -2739 1315
rect -2811 1261 -2739 1281
rect -2465 1315 -2393 1481
rect -2465 1281 -2451 1315
rect -2417 1281 -2393 1315
rect -2465 1261 -2393 1281
rect -2811 1247 -2393 1261
rect -2811 1213 -2787 1247
rect -2753 1213 -2719 1247
rect -2685 1213 -2519 1247
rect -2485 1213 -2451 1247
rect -2417 1213 -2393 1247
rect -2811 1189 -2393 1213
rect -2331 1600 -2230 1634
rect -2331 1566 -2298 1600
rect -2264 1566 -2230 1600
rect -2331 1532 -2230 1566
rect -2331 1498 -2298 1532
rect -2264 1498 -2230 1532
rect -2331 1298 -2230 1498
rect -2331 1264 -2298 1298
rect -2264 1264 -2230 1298
rect -2331 1230 -2230 1264
rect -2331 1196 -2298 1230
rect -2264 1196 -2230 1230
rect -2974 1128 -2940 1162
rect -2906 1128 -2873 1162
rect -2974 1127 -2873 1128
rect -2331 1162 -2230 1196
rect -2331 1128 -2298 1162
rect -2264 1128 -2230 1162
rect -2331 1127 -2230 1128
rect -2974 1094 -2230 1127
rect -2974 1060 -2940 1094
rect -2906 1060 -2872 1094
rect -2838 1060 -2804 1094
rect -2770 1060 -2736 1094
rect -2702 1060 -2502 1094
rect -2468 1060 -2434 1094
rect -2400 1060 -2366 1094
rect -2332 1060 -2298 1094
rect -2264 1060 -2230 1094
rect -2974 1026 -2230 1060
rect -1974 1736 -1230 1770
rect -1974 1702 -1940 1736
rect -1906 1702 -1872 1736
rect -1838 1702 -1804 1736
rect -1770 1702 -1736 1736
rect -1702 1702 -1502 1736
rect -1468 1702 -1434 1736
rect -1400 1702 -1366 1736
rect -1332 1702 -1298 1736
rect -1264 1702 -1230 1736
rect -1974 1669 -1230 1702
rect -1974 1668 -1873 1669
rect -1974 1634 -1940 1668
rect -1906 1634 -1873 1668
rect -1974 1600 -1873 1634
rect -1331 1668 -1230 1669
rect -1331 1634 -1298 1668
rect -1264 1634 -1230 1668
rect -1974 1566 -1940 1600
rect -1906 1566 -1873 1600
rect -1974 1532 -1873 1566
rect -1974 1498 -1940 1532
rect -1906 1498 -1873 1532
rect -1974 1298 -1873 1498
rect -1974 1264 -1940 1298
rect -1906 1264 -1873 1298
rect -1974 1230 -1873 1264
rect -1974 1196 -1940 1230
rect -1906 1196 -1873 1230
rect -1974 1162 -1873 1196
rect -1811 1583 -1393 1607
rect -1811 1549 -1787 1583
rect -1753 1549 -1719 1583
rect -1685 1549 -1519 1583
rect -1485 1549 -1451 1583
rect -1417 1549 -1393 1583
rect -1811 1535 -1393 1549
rect -1811 1515 -1739 1535
rect -1811 1481 -1787 1515
rect -1753 1481 -1739 1515
rect -1811 1315 -1739 1481
rect -1465 1515 -1393 1535
rect -1465 1481 -1451 1515
rect -1417 1481 -1393 1515
rect -1681 1463 -1523 1477
rect -1681 1429 -1667 1463
rect -1633 1449 -1571 1463
rect -1537 1429 -1523 1463
rect -1681 1367 -1653 1429
rect -1551 1367 -1523 1429
rect -1681 1333 -1667 1367
rect -1633 1333 -1571 1347
rect -1537 1333 -1523 1367
rect -1681 1319 -1523 1333
rect -1811 1281 -1787 1315
rect -1753 1281 -1739 1315
rect -1811 1261 -1739 1281
rect -1465 1315 -1393 1481
rect -1465 1281 -1451 1315
rect -1417 1281 -1393 1315
rect -1465 1261 -1393 1281
rect -1811 1247 -1393 1261
rect -1811 1213 -1787 1247
rect -1753 1213 -1719 1247
rect -1685 1213 -1519 1247
rect -1485 1213 -1451 1247
rect -1417 1213 -1393 1247
rect -1811 1189 -1393 1213
rect -1331 1600 -1230 1634
rect -1331 1566 -1298 1600
rect -1264 1566 -1230 1600
rect -1331 1532 -1230 1566
rect -1331 1498 -1298 1532
rect -1264 1498 -1230 1532
rect -1331 1298 -1230 1498
rect -1331 1264 -1298 1298
rect -1264 1264 -1230 1298
rect -1331 1230 -1230 1264
rect -1331 1196 -1298 1230
rect -1264 1196 -1230 1230
rect -1974 1128 -1940 1162
rect -1906 1128 -1873 1162
rect -1974 1127 -1873 1128
rect -1331 1162 -1230 1196
rect -1331 1128 -1298 1162
rect -1264 1128 -1230 1162
rect -1331 1127 -1230 1128
rect -1974 1094 -1230 1127
rect -1974 1060 -1940 1094
rect -1906 1060 -1872 1094
rect -1838 1060 -1804 1094
rect -1770 1060 -1736 1094
rect -1702 1060 -1502 1094
rect -1468 1060 -1434 1094
rect -1400 1060 -1366 1094
rect -1332 1060 -1298 1094
rect -1264 1060 -1230 1094
rect -1974 1026 -1230 1060
rect -974 1736 -230 1770
rect -974 1702 -940 1736
rect -906 1702 -872 1736
rect -838 1702 -804 1736
rect -770 1702 -736 1736
rect -702 1702 -502 1736
rect -468 1702 -434 1736
rect -400 1702 -366 1736
rect -332 1702 -298 1736
rect -264 1702 -230 1736
rect -974 1669 -230 1702
rect -974 1668 -873 1669
rect -974 1634 -940 1668
rect -906 1634 -873 1668
rect -974 1600 -873 1634
rect -331 1668 -230 1669
rect -331 1634 -298 1668
rect -264 1634 -230 1668
rect -974 1566 -940 1600
rect -906 1566 -873 1600
rect -974 1532 -873 1566
rect -974 1498 -940 1532
rect -906 1498 -873 1532
rect -974 1298 -873 1498
rect -974 1264 -940 1298
rect -906 1264 -873 1298
rect -974 1230 -873 1264
rect -974 1196 -940 1230
rect -906 1196 -873 1230
rect -974 1162 -873 1196
rect -811 1583 -393 1607
rect -811 1549 -787 1583
rect -753 1549 -719 1583
rect -685 1549 -519 1583
rect -485 1549 -451 1583
rect -417 1549 -393 1583
rect -811 1535 -393 1549
rect -811 1515 -739 1535
rect -811 1481 -787 1515
rect -753 1481 -739 1515
rect -811 1315 -739 1481
rect -465 1515 -393 1535
rect -465 1481 -451 1515
rect -417 1481 -393 1515
rect -681 1463 -523 1477
rect -681 1429 -667 1463
rect -633 1449 -571 1463
rect -537 1429 -523 1463
rect -681 1367 -653 1429
rect -551 1367 -523 1429
rect -681 1333 -667 1367
rect -633 1333 -571 1347
rect -537 1333 -523 1367
rect -681 1319 -523 1333
rect -811 1281 -787 1315
rect -753 1281 -739 1315
rect -811 1261 -739 1281
rect -465 1315 -393 1481
rect -465 1281 -451 1315
rect -417 1281 -393 1315
rect -465 1261 -393 1281
rect -811 1247 -393 1261
rect -811 1213 -787 1247
rect -753 1213 -719 1247
rect -685 1213 -519 1247
rect -485 1213 -451 1247
rect -417 1213 -393 1247
rect -811 1189 -393 1213
rect -331 1600 -230 1634
rect -331 1566 -298 1600
rect -264 1566 -230 1600
rect -331 1532 -230 1566
rect -331 1498 -298 1532
rect -264 1498 -230 1532
rect -331 1298 -230 1498
rect -331 1264 -298 1298
rect -264 1264 -230 1298
rect -331 1230 -230 1264
rect -331 1196 -298 1230
rect -264 1196 -230 1230
rect -974 1128 -940 1162
rect -906 1128 -873 1162
rect -974 1127 -873 1128
rect -331 1162 -230 1196
rect -331 1128 -298 1162
rect -264 1128 -230 1162
rect -331 1127 -230 1128
rect -974 1094 -230 1127
rect -974 1060 -940 1094
rect -906 1060 -872 1094
rect -838 1060 -804 1094
rect -770 1060 -736 1094
rect -702 1060 -502 1094
rect -468 1060 -434 1094
rect -400 1060 -366 1094
rect -332 1060 -298 1094
rect -264 1060 -230 1094
rect -974 1026 -230 1060
rect 26 1736 770 1770
rect 26 1702 60 1736
rect 94 1702 128 1736
rect 162 1702 196 1736
rect 230 1702 264 1736
rect 298 1702 498 1736
rect 532 1702 566 1736
rect 600 1702 634 1736
rect 668 1702 702 1736
rect 736 1702 770 1736
rect 26 1669 770 1702
rect 26 1668 127 1669
rect 26 1634 60 1668
rect 94 1634 127 1668
rect 26 1600 127 1634
rect 669 1668 770 1669
rect 669 1634 702 1668
rect 736 1634 770 1668
rect 26 1566 60 1600
rect 94 1566 127 1600
rect 26 1532 127 1566
rect 26 1498 60 1532
rect 94 1498 127 1532
rect 26 1298 127 1498
rect 26 1264 60 1298
rect 94 1264 127 1298
rect 26 1230 127 1264
rect 26 1196 60 1230
rect 94 1196 127 1230
rect 26 1162 127 1196
rect 189 1583 607 1607
rect 189 1549 213 1583
rect 247 1549 281 1583
rect 315 1549 481 1583
rect 515 1549 549 1583
rect 583 1549 607 1583
rect 189 1535 607 1549
rect 189 1515 261 1535
rect 189 1481 213 1515
rect 247 1481 261 1515
rect 189 1315 261 1481
rect 535 1515 607 1535
rect 535 1481 549 1515
rect 583 1481 607 1515
rect 319 1463 477 1477
rect 319 1429 333 1463
rect 367 1449 429 1463
rect 463 1429 477 1463
rect 319 1367 347 1429
rect 449 1367 477 1429
rect 319 1333 333 1367
rect 367 1333 429 1347
rect 463 1333 477 1367
rect 319 1319 477 1333
rect 189 1281 213 1315
rect 247 1281 261 1315
rect 189 1261 261 1281
rect 535 1315 607 1481
rect 535 1281 549 1315
rect 583 1281 607 1315
rect 535 1261 607 1281
rect 189 1247 607 1261
rect 189 1213 213 1247
rect 247 1213 281 1247
rect 315 1213 481 1247
rect 515 1213 549 1247
rect 583 1213 607 1247
rect 189 1189 607 1213
rect 669 1600 770 1634
rect 669 1566 702 1600
rect 736 1566 770 1600
rect 669 1532 770 1566
rect 669 1498 702 1532
rect 736 1498 770 1532
rect 669 1298 770 1498
rect 669 1264 702 1298
rect 736 1264 770 1298
rect 669 1230 770 1264
rect 669 1196 702 1230
rect 736 1196 770 1230
rect 26 1128 60 1162
rect 94 1128 127 1162
rect 26 1127 127 1128
rect 669 1162 770 1196
rect 669 1128 702 1162
rect 736 1128 770 1162
rect 669 1127 770 1128
rect 26 1094 770 1127
rect 26 1060 60 1094
rect 94 1060 128 1094
rect 162 1060 196 1094
rect 230 1060 264 1094
rect 298 1060 498 1094
rect 532 1060 566 1094
rect 600 1060 634 1094
rect 668 1060 702 1094
rect 736 1060 770 1094
rect 26 1026 770 1060
rect 1026 1736 1770 1770
rect 1026 1702 1060 1736
rect 1094 1702 1128 1736
rect 1162 1702 1196 1736
rect 1230 1702 1264 1736
rect 1298 1702 1498 1736
rect 1532 1702 1566 1736
rect 1600 1702 1634 1736
rect 1668 1702 1702 1736
rect 1736 1702 1770 1736
rect 1026 1669 1770 1702
rect 1026 1668 1127 1669
rect 1026 1634 1060 1668
rect 1094 1634 1127 1668
rect 1026 1600 1127 1634
rect 1669 1668 1770 1669
rect 1669 1634 1702 1668
rect 1736 1634 1770 1668
rect 1026 1566 1060 1600
rect 1094 1566 1127 1600
rect 1026 1532 1127 1566
rect 1026 1498 1060 1532
rect 1094 1498 1127 1532
rect 1026 1298 1127 1498
rect 1026 1264 1060 1298
rect 1094 1264 1127 1298
rect 1026 1230 1127 1264
rect 1026 1196 1060 1230
rect 1094 1196 1127 1230
rect 1026 1162 1127 1196
rect 1189 1583 1607 1607
rect 1189 1549 1213 1583
rect 1247 1549 1281 1583
rect 1315 1549 1481 1583
rect 1515 1549 1549 1583
rect 1583 1549 1607 1583
rect 1189 1535 1607 1549
rect 1189 1515 1261 1535
rect 1189 1481 1213 1515
rect 1247 1481 1261 1515
rect 1189 1315 1261 1481
rect 1535 1515 1607 1535
rect 1535 1481 1549 1515
rect 1583 1481 1607 1515
rect 1319 1463 1477 1477
rect 1319 1429 1333 1463
rect 1367 1449 1429 1463
rect 1463 1429 1477 1463
rect 1319 1367 1347 1429
rect 1449 1367 1477 1429
rect 1319 1333 1333 1367
rect 1367 1333 1429 1347
rect 1463 1333 1477 1367
rect 1319 1319 1477 1333
rect 1189 1281 1213 1315
rect 1247 1281 1261 1315
rect 1189 1261 1261 1281
rect 1535 1315 1607 1481
rect 1535 1281 1549 1315
rect 1583 1281 1607 1315
rect 1535 1261 1607 1281
rect 1189 1247 1607 1261
rect 1189 1213 1213 1247
rect 1247 1213 1281 1247
rect 1315 1213 1481 1247
rect 1515 1213 1549 1247
rect 1583 1213 1607 1247
rect 1189 1189 1607 1213
rect 1669 1600 1770 1634
rect 1669 1566 1702 1600
rect 1736 1566 1770 1600
rect 1669 1532 1770 1566
rect 1669 1498 1702 1532
rect 1736 1498 1770 1532
rect 1669 1298 1770 1498
rect 1669 1264 1702 1298
rect 1736 1264 1770 1298
rect 1669 1230 1770 1264
rect 1669 1196 1702 1230
rect 1736 1196 1770 1230
rect 1026 1128 1060 1162
rect 1094 1128 1127 1162
rect 1026 1127 1127 1128
rect 1669 1162 1770 1196
rect 1669 1128 1702 1162
rect 1736 1128 1770 1162
rect 1669 1127 1770 1128
rect 1026 1094 1770 1127
rect 1026 1060 1060 1094
rect 1094 1060 1128 1094
rect 1162 1060 1196 1094
rect 1230 1060 1264 1094
rect 1298 1060 1498 1094
rect 1532 1060 1566 1094
rect 1600 1060 1634 1094
rect 1668 1060 1702 1094
rect 1736 1060 1770 1094
rect 1026 1026 1770 1060
rect -3974 736 -3230 770
rect -3974 702 -3940 736
rect -3906 702 -3872 736
rect -3838 702 -3804 736
rect -3770 702 -3736 736
rect -3702 702 -3502 736
rect -3468 702 -3434 736
rect -3400 702 -3366 736
rect -3332 702 -3298 736
rect -3264 702 -3230 736
rect -3974 669 -3230 702
rect -3974 668 -3873 669
rect -3974 634 -3940 668
rect -3906 634 -3873 668
rect -3974 600 -3873 634
rect -3331 668 -3230 669
rect -3331 634 -3298 668
rect -3264 634 -3230 668
rect -3974 566 -3940 600
rect -3906 566 -3873 600
rect -3974 532 -3873 566
rect -3974 498 -3940 532
rect -3906 498 -3873 532
rect -3974 298 -3873 498
rect -3974 264 -3940 298
rect -3906 264 -3873 298
rect -3974 230 -3873 264
rect -3974 196 -3940 230
rect -3906 196 -3873 230
rect -3974 162 -3873 196
rect -3811 583 -3393 607
rect -3811 549 -3787 583
rect -3753 549 -3719 583
rect -3685 549 -3519 583
rect -3485 549 -3451 583
rect -3417 549 -3393 583
rect -3811 535 -3393 549
rect -3811 515 -3739 535
rect -3811 481 -3787 515
rect -3753 481 -3739 515
rect -3811 315 -3739 481
rect -3465 515 -3393 535
rect -3465 481 -3451 515
rect -3417 481 -3393 515
rect -3681 463 -3523 477
rect -3681 429 -3667 463
rect -3633 449 -3571 463
rect -3537 429 -3523 463
rect -3681 367 -3653 429
rect -3551 367 -3523 429
rect -3681 333 -3667 367
rect -3633 333 -3571 347
rect -3537 333 -3523 367
rect -3681 319 -3523 333
rect -3811 281 -3787 315
rect -3753 281 -3739 315
rect -3811 261 -3739 281
rect -3465 315 -3393 481
rect -3465 281 -3451 315
rect -3417 281 -3393 315
rect -3465 261 -3393 281
rect -3811 247 -3393 261
rect -3811 213 -3787 247
rect -3753 213 -3719 247
rect -3685 213 -3519 247
rect -3485 213 -3451 247
rect -3417 213 -3393 247
rect -3811 189 -3393 213
rect -3331 600 -3230 634
rect -3331 566 -3298 600
rect -3264 566 -3230 600
rect -3331 532 -3230 566
rect -3331 498 -3298 532
rect -3264 498 -3230 532
rect -3331 298 -3230 498
rect -3331 264 -3298 298
rect -3264 264 -3230 298
rect -3331 230 -3230 264
rect -3331 196 -3298 230
rect -3264 196 -3230 230
rect -3974 128 -3940 162
rect -3906 128 -3873 162
rect -3974 127 -3873 128
rect -3331 162 -3230 196
rect -3331 128 -3298 162
rect -3264 128 -3230 162
rect -3331 127 -3230 128
rect -3974 94 -3230 127
rect -3974 60 -3940 94
rect -3906 60 -3872 94
rect -3838 60 -3804 94
rect -3770 60 -3736 94
rect -3702 60 -3502 94
rect -3468 60 -3434 94
rect -3400 60 -3366 94
rect -3332 60 -3298 94
rect -3264 60 -3230 94
rect -3974 26 -3230 60
rect -2974 736 -230 770
rect -2974 702 -2940 736
rect -2906 702 -2872 736
rect -2838 702 -2804 736
rect -2770 702 -2736 736
rect -2702 702 -2502 736
rect -2468 702 -2434 736
rect -2400 702 -2366 736
rect -2332 702 -2298 736
rect -2264 702 -1940 736
rect -1906 702 -1872 736
rect -1838 702 -1804 736
rect -1770 702 -1736 736
rect -1702 702 -1502 736
rect -1468 702 -1434 736
rect -1400 702 -1366 736
rect -1332 702 -1298 736
rect -1264 702 -940 736
rect -906 702 -872 736
rect -838 702 -804 736
rect -770 702 -736 736
rect -702 702 -502 736
rect -468 702 -434 736
rect -400 702 -366 736
rect -332 702 -298 736
rect -264 702 -230 736
rect -2974 670 -230 702
rect -2974 669 -2230 670
rect -2974 668 -2873 669
rect -2974 634 -2940 668
rect -2906 634 -2873 668
rect -2974 600 -2873 634
rect -2331 668 -2230 669
rect -2331 634 -2298 668
rect -2264 634 -2230 668
rect -2331 610 -2230 634
rect -2120 610 -2080 670
rect -1974 669 -1230 670
rect -1974 668 -1873 669
rect -1974 634 -1940 668
rect -1906 634 -1873 668
rect -1974 610 -1873 634
rect -1331 668 -1230 669
rect -1331 634 -1298 668
rect -1264 634 -1230 668
rect -1331 610 -1230 634
rect -1120 610 -1080 670
rect -974 669 -230 670
rect -974 668 -873 669
rect -974 634 -940 668
rect -906 634 -873 668
rect -974 610 -873 634
rect -331 668 -230 669
rect -331 634 -298 668
rect -264 634 -230 668
rect -2490 607 -770 610
rect -2974 566 -2940 600
rect -2906 566 -2873 600
rect -2974 532 -2873 566
rect -2974 498 -2940 532
rect -2906 498 -2873 532
rect -2974 298 -2873 498
rect -2974 264 -2940 298
rect -2906 264 -2873 298
rect -2974 230 -2873 264
rect -2974 196 -2940 230
rect -2906 196 -2873 230
rect -2974 162 -2873 196
rect -2811 600 -393 607
rect -2811 583 -2298 600
rect -2811 549 -2787 583
rect -2753 549 -2719 583
rect -2685 549 -2519 583
rect -2485 549 -2451 583
rect -2417 566 -2298 583
rect -2264 566 -1940 600
rect -1906 583 -1298 600
rect -1906 566 -1787 583
rect -2417 549 -1787 566
rect -1753 549 -1719 583
rect -1685 549 -1519 583
rect -1485 549 -1451 583
rect -1417 566 -1298 583
rect -1264 566 -940 600
rect -906 583 -393 600
rect -906 566 -787 583
rect -1417 549 -787 566
rect -753 549 -719 583
rect -685 549 -519 583
rect -485 549 -451 583
rect -417 549 -393 583
rect -2811 535 -393 549
rect -2811 515 -2739 535
rect -2490 532 -739 535
rect -2490 530 -2298 532
rect -2811 481 -2787 515
rect -2753 481 -2739 515
rect -2811 315 -2739 481
rect -2465 515 -2393 530
rect -2465 481 -2451 515
rect -2417 481 -2393 515
rect -2681 463 -2523 477
rect -2681 429 -2667 463
rect -2633 449 -2571 463
rect -2537 429 -2523 463
rect -2681 367 -2653 429
rect -2551 367 -2523 429
rect -2681 333 -2667 367
rect -2633 333 -2571 347
rect -2537 333 -2523 367
rect -2681 319 -2523 333
rect -2811 281 -2787 315
rect -2753 281 -2739 315
rect -2811 261 -2739 281
rect -2465 315 -2393 481
rect -2465 281 -2451 315
rect -2417 281 -2393 315
rect -2465 261 -2393 281
rect -2811 247 -2393 261
rect -2811 213 -2787 247
rect -2753 213 -2719 247
rect -2685 213 -2519 247
rect -2485 213 -2451 247
rect -2417 213 -2393 247
rect -2811 189 -2393 213
rect -2331 498 -2298 530
rect -2264 530 -1940 532
rect -2264 498 -2230 530
rect -2331 298 -2230 498
rect -2331 264 -2298 298
rect -2264 264 -2230 298
rect -2331 230 -2230 264
rect -2331 196 -2298 230
rect -2264 196 -2230 230
rect -2974 128 -2940 162
rect -2906 128 -2873 162
rect -2974 127 -2873 128
rect -2331 162 -2230 196
rect -2331 128 -2298 162
rect -2264 128 -2230 162
rect -2331 127 -2230 128
rect -2974 94 -2230 127
rect -2974 60 -2940 94
rect -2906 60 -2872 94
rect -2838 60 -2804 94
rect -2770 60 -2736 94
rect -2702 60 -2502 94
rect -2468 60 -2434 94
rect -2400 60 -2366 94
rect -2332 60 -2298 94
rect -2264 60 -2230 94
rect -2974 26 -2230 60
rect -2120 -230 -2080 530
rect -1974 498 -1940 530
rect -1906 530 -1298 532
rect -1906 498 -1873 530
rect -1974 298 -1873 498
rect -1974 264 -1940 298
rect -1906 264 -1873 298
rect -1974 230 -1873 264
rect -1974 196 -1940 230
rect -1906 196 -1873 230
rect -1974 162 -1873 196
rect -1811 515 -1739 530
rect -1811 481 -1787 515
rect -1753 481 -1739 515
rect -1811 315 -1739 481
rect -1465 515 -1393 530
rect -1465 481 -1451 515
rect -1417 481 -1393 515
rect -1681 463 -1523 477
rect -1681 429 -1667 463
rect -1633 449 -1571 463
rect -1537 429 -1523 463
rect -1681 367 -1653 429
rect -1551 367 -1523 429
rect -1681 333 -1667 367
rect -1633 333 -1571 347
rect -1537 333 -1523 367
rect -1681 319 -1523 333
rect -1811 281 -1787 315
rect -1753 281 -1739 315
rect -1811 261 -1739 281
rect -1465 315 -1393 481
rect -1465 281 -1451 315
rect -1417 281 -1393 315
rect -1465 261 -1393 281
rect -1811 247 -1393 261
rect -1811 213 -1787 247
rect -1753 213 -1719 247
rect -1685 213 -1519 247
rect -1485 213 -1451 247
rect -1417 213 -1393 247
rect -1811 189 -1393 213
rect -1331 498 -1298 530
rect -1264 530 -940 532
rect -1264 498 -1230 530
rect -1331 298 -1230 498
rect -1331 264 -1298 298
rect -1264 264 -1230 298
rect -1331 230 -1230 264
rect -1331 196 -1298 230
rect -1264 196 -1230 230
rect -1974 128 -1940 162
rect -1906 128 -1873 162
rect -1974 127 -1873 128
rect -1331 162 -1230 196
rect -1331 128 -1298 162
rect -1264 128 -1230 162
rect -1331 127 -1230 128
rect -1974 94 -1230 127
rect -1974 60 -1940 94
rect -1906 60 -1872 94
rect -1838 60 -1804 94
rect -1770 60 -1736 94
rect -1702 60 -1502 94
rect -1468 60 -1434 94
rect -1400 60 -1366 94
rect -1332 60 -1298 94
rect -1264 60 -1230 94
rect -1974 26 -1230 60
rect -1120 -230 -1080 530
rect -974 498 -940 530
rect -906 530 -739 532
rect -906 498 -873 530
rect -974 298 -873 498
rect -974 264 -940 298
rect -906 264 -873 298
rect -974 230 -873 264
rect -974 196 -940 230
rect -906 196 -873 230
rect -974 162 -873 196
rect -811 515 -739 530
rect -811 481 -787 515
rect -753 481 -739 515
rect -811 315 -739 481
rect -465 515 -393 535
rect -465 481 -451 515
rect -417 481 -393 515
rect -681 463 -523 477
rect -681 429 -667 463
rect -633 449 -571 463
rect -537 429 -523 463
rect -681 367 -653 429
rect -551 367 -523 429
rect -681 333 -667 367
rect -633 333 -571 347
rect -537 333 -523 367
rect -681 319 -523 333
rect -811 281 -787 315
rect -753 281 -739 315
rect -811 261 -739 281
rect -465 315 -393 481
rect -465 281 -451 315
rect -417 281 -393 315
rect -465 261 -393 281
rect -811 247 -393 261
rect -811 213 -787 247
rect -753 213 -719 247
rect -685 213 -519 247
rect -485 213 -451 247
rect -417 213 -393 247
rect -811 189 -393 213
rect -331 600 -230 634
rect -331 566 -298 600
rect -264 566 -230 600
rect -331 532 -230 566
rect -331 498 -298 532
rect -264 498 -230 532
rect -331 298 -230 498
rect -331 264 -298 298
rect -264 264 -230 298
rect -331 230 -230 264
rect -331 196 -298 230
rect -264 196 -230 230
rect -974 128 -940 162
rect -906 128 -873 162
rect -974 127 -873 128
rect -331 162 -230 196
rect -331 128 -298 162
rect -264 128 -230 162
rect -331 127 -230 128
rect -974 94 -230 127
rect -974 60 -940 94
rect -906 60 -872 94
rect -838 60 -804 94
rect -770 60 -736 94
rect -702 60 -502 94
rect -468 60 -434 94
rect -400 60 -366 94
rect -332 60 -298 94
rect -264 60 -230 94
rect -974 26 -230 60
rect 26 736 770 770
rect 26 702 60 736
rect 94 702 128 736
rect 162 702 196 736
rect 230 702 264 736
rect 298 702 498 736
rect 532 702 566 736
rect 600 702 634 736
rect 668 702 702 736
rect 736 702 770 736
rect 26 669 770 702
rect 26 668 127 669
rect 26 634 60 668
rect 94 634 127 668
rect 26 600 127 634
rect 669 668 770 669
rect 669 634 702 668
rect 736 634 770 668
rect 26 566 60 600
rect 94 566 127 600
rect 26 532 127 566
rect 26 498 60 532
rect 94 498 127 532
rect 26 298 127 498
rect 26 264 60 298
rect 94 264 127 298
rect 26 230 127 264
rect 26 196 60 230
rect 94 196 127 230
rect 26 162 127 196
rect 189 583 607 607
rect 189 549 213 583
rect 247 549 281 583
rect 315 549 481 583
rect 515 549 549 583
rect 583 549 607 583
rect 189 535 607 549
rect 189 515 261 535
rect 189 481 213 515
rect 247 481 261 515
rect 189 315 261 481
rect 535 515 607 535
rect 535 481 549 515
rect 583 481 607 515
rect 319 463 477 477
rect 319 429 333 463
rect 367 449 429 463
rect 463 429 477 463
rect 319 367 347 429
rect 449 367 477 429
rect 319 333 333 367
rect 367 333 429 347
rect 463 333 477 367
rect 319 319 477 333
rect 189 281 213 315
rect 247 281 261 315
rect 189 261 261 281
rect 535 315 607 481
rect 535 281 549 315
rect 583 281 607 315
rect 535 261 607 281
rect 189 247 607 261
rect 189 213 213 247
rect 247 213 281 247
rect 315 213 481 247
rect 515 213 549 247
rect 583 213 607 247
rect 189 189 607 213
rect 669 600 770 634
rect 669 566 702 600
rect 736 566 770 600
rect 669 532 770 566
rect 669 498 702 532
rect 736 498 770 532
rect 669 298 770 498
rect 669 264 702 298
rect 736 264 770 298
rect 669 230 770 264
rect 669 196 702 230
rect 736 196 770 230
rect 26 128 60 162
rect 94 128 127 162
rect 26 127 127 128
rect 669 162 770 196
rect 669 128 702 162
rect 736 128 770 162
rect 669 127 770 128
rect 26 94 770 127
rect 26 60 60 94
rect 94 60 128 94
rect 162 60 196 94
rect 230 60 264 94
rect 298 60 498 94
rect 532 60 566 94
rect 600 60 634 94
rect 668 60 702 94
rect 736 60 770 94
rect 26 26 770 60
rect 1026 736 1770 770
rect 1026 702 1060 736
rect 1094 702 1128 736
rect 1162 702 1196 736
rect 1230 702 1264 736
rect 1298 702 1498 736
rect 1532 702 1566 736
rect 1600 702 1634 736
rect 1668 702 1702 736
rect 1736 702 1770 736
rect 1026 669 1770 702
rect 1026 668 1127 669
rect 1026 634 1060 668
rect 1094 634 1127 668
rect 1026 600 1127 634
rect 1669 668 1770 669
rect 1669 634 1702 668
rect 1736 634 1770 668
rect 1026 566 1060 600
rect 1094 566 1127 600
rect 1026 532 1127 566
rect 1026 498 1060 532
rect 1094 498 1127 532
rect 1026 298 1127 498
rect 1026 264 1060 298
rect 1094 264 1127 298
rect 1026 230 1127 264
rect 1026 196 1060 230
rect 1094 196 1127 230
rect 1026 162 1127 196
rect 1189 583 1607 607
rect 1189 549 1213 583
rect 1247 549 1281 583
rect 1315 549 1481 583
rect 1515 549 1549 583
rect 1583 549 1607 583
rect 1189 535 1607 549
rect 1189 515 1261 535
rect 1189 481 1213 515
rect 1247 481 1261 515
rect 1189 315 1261 481
rect 1535 515 1607 535
rect 1535 481 1549 515
rect 1583 481 1607 515
rect 1319 463 1477 477
rect 1319 429 1333 463
rect 1367 449 1429 463
rect 1463 429 1477 463
rect 1319 367 1347 429
rect 1449 367 1477 429
rect 1319 333 1333 367
rect 1367 333 1429 347
rect 1463 333 1477 367
rect 1319 319 1477 333
rect 1189 281 1213 315
rect 1247 281 1261 315
rect 1189 261 1261 281
rect 1535 315 1607 481
rect 1535 281 1549 315
rect 1583 281 1607 315
rect 1535 261 1607 281
rect 1189 247 1607 261
rect 1189 213 1213 247
rect 1247 213 1281 247
rect 1315 213 1481 247
rect 1515 213 1549 247
rect 1583 213 1607 247
rect 1189 189 1607 213
rect 1669 600 1770 634
rect 1669 566 1702 600
rect 1736 566 1770 600
rect 1669 532 1770 566
rect 1669 498 1702 532
rect 1736 498 1770 532
rect 1669 298 1770 498
rect 1669 264 1702 298
rect 1736 264 1770 298
rect 1669 230 1770 264
rect 1669 196 1702 230
rect 1736 196 1770 230
rect 1026 128 1060 162
rect 1094 128 1127 162
rect 1026 127 1127 128
rect 1669 162 1770 196
rect 1669 128 1702 162
rect 1736 128 1770 162
rect 1669 127 1770 128
rect 1026 94 1770 127
rect 1026 60 1060 94
rect 1094 60 1128 94
rect 1162 60 1196 94
rect 1230 60 1264 94
rect 1298 60 1498 94
rect 1532 60 1566 94
rect 1600 60 1634 94
rect 1668 60 1702 94
rect 1736 60 1770 94
rect 1026 26 1770 60
rect -3974 -264 -3230 -230
rect -3974 -298 -3940 -264
rect -3906 -298 -3872 -264
rect -3838 -298 -3804 -264
rect -3770 -298 -3736 -264
rect -3702 -298 -3502 -264
rect -3468 -298 -3434 -264
rect -3400 -298 -3366 -264
rect -3332 -298 -3298 -264
rect -3264 -298 -3230 -264
rect -3974 -331 -3230 -298
rect -3974 -332 -3873 -331
rect -3974 -366 -3940 -332
rect -3906 -366 -3873 -332
rect -3974 -400 -3873 -366
rect -3331 -332 -3230 -331
rect -3331 -366 -3298 -332
rect -3264 -366 -3230 -332
rect -3974 -434 -3940 -400
rect -3906 -434 -3873 -400
rect -3974 -468 -3873 -434
rect -3974 -502 -3940 -468
rect -3906 -502 -3873 -468
rect -3974 -702 -3873 -502
rect -3974 -736 -3940 -702
rect -3906 -736 -3873 -702
rect -3974 -770 -3873 -736
rect -3974 -804 -3940 -770
rect -3906 -804 -3873 -770
rect -3974 -838 -3873 -804
rect -3811 -417 -3393 -393
rect -3811 -451 -3787 -417
rect -3753 -451 -3719 -417
rect -3685 -451 -3519 -417
rect -3485 -451 -3451 -417
rect -3417 -451 -3393 -417
rect -3811 -465 -3393 -451
rect -3811 -485 -3739 -465
rect -3811 -519 -3787 -485
rect -3753 -519 -3739 -485
rect -3811 -685 -3739 -519
rect -3465 -485 -3393 -465
rect -3465 -519 -3451 -485
rect -3417 -519 -3393 -485
rect -3681 -537 -3523 -523
rect -3681 -571 -3667 -537
rect -3633 -551 -3571 -537
rect -3537 -571 -3523 -537
rect -3681 -633 -3653 -571
rect -3551 -633 -3523 -571
rect -3681 -667 -3667 -633
rect -3633 -667 -3571 -653
rect -3537 -667 -3523 -633
rect -3681 -681 -3523 -667
rect -3811 -719 -3787 -685
rect -3753 -719 -3739 -685
rect -3811 -739 -3739 -719
rect -3465 -685 -3393 -519
rect -3465 -719 -3451 -685
rect -3417 -719 -3393 -685
rect -3465 -739 -3393 -719
rect -3811 -753 -3393 -739
rect -3811 -787 -3787 -753
rect -3753 -787 -3719 -753
rect -3685 -787 -3519 -753
rect -3485 -787 -3451 -753
rect -3417 -787 -3393 -753
rect -3811 -811 -3393 -787
rect -3331 -400 -3230 -366
rect -3331 -434 -3298 -400
rect -3264 -434 -3230 -400
rect -3331 -468 -3230 -434
rect -3331 -502 -3298 -468
rect -3264 -502 -3230 -468
rect -3331 -702 -3230 -502
rect -3331 -736 -3298 -702
rect -3264 -736 -3230 -702
rect -3331 -770 -3230 -736
rect -3331 -804 -3298 -770
rect -3264 -804 -3230 -770
rect -3974 -872 -3940 -838
rect -3906 -872 -3873 -838
rect -3974 -873 -3873 -872
rect -3331 -838 -3230 -804
rect -3331 -872 -3298 -838
rect -3264 -872 -3230 -838
rect -3331 -873 -3230 -872
rect -3974 -906 -3230 -873
rect -3974 -940 -3940 -906
rect -3906 -940 -3872 -906
rect -3838 -940 -3804 -906
rect -3770 -940 -3736 -906
rect -3702 -940 -3502 -906
rect -3468 -940 -3434 -906
rect -3400 -940 -3366 -906
rect -3332 -940 -3298 -906
rect -3264 -940 -3230 -906
rect -3974 -974 -3230 -940
rect -2974 -264 -230 -230
rect -2974 -298 -2940 -264
rect -2906 -298 -2872 -264
rect -2838 -298 -2804 -264
rect -2770 -298 -2736 -264
rect -2702 -298 -2502 -264
rect -2468 -298 -2434 -264
rect -2400 -298 -2366 -264
rect -2332 -298 -2298 -264
rect -2264 -298 -1940 -264
rect -1906 -298 -1872 -264
rect -1838 -298 -1804 -264
rect -1770 -298 -1736 -264
rect -1702 -298 -1502 -264
rect -1468 -298 -1434 -264
rect -1400 -298 -1366 -264
rect -1332 -298 -1298 -264
rect -1264 -298 -940 -264
rect -906 -298 -872 -264
rect -838 -298 -804 -264
rect -770 -298 -736 -264
rect -702 -298 -502 -264
rect -468 -298 -434 -264
rect -400 -298 -366 -264
rect -332 -298 -298 -264
rect -264 -298 -230 -264
rect -2974 -331 -230 -298
rect -2974 -332 -2873 -331
rect -2974 -366 -2940 -332
rect -2906 -366 -2873 -332
rect -2390 -332 -750 -331
rect -2390 -340 -2298 -332
rect -2974 -400 -2873 -366
rect -2331 -366 -2298 -340
rect -2264 -340 -1940 -332
rect -2264 -366 -2230 -340
rect -2331 -390 -2230 -366
rect -2120 -390 -2080 -340
rect -1974 -366 -1940 -340
rect -1906 -340 -1298 -332
rect -1906 -366 -1873 -340
rect -1974 -390 -1873 -366
rect -1331 -366 -1298 -340
rect -1264 -340 -940 -332
rect -1264 -366 -1230 -340
rect -1331 -390 -1230 -366
rect -1120 -390 -1080 -340
rect -974 -366 -940 -340
rect -906 -340 -750 -332
rect -331 -332 -230 -331
rect -906 -366 -873 -340
rect -974 -390 -873 -366
rect -331 -366 -298 -332
rect -264 -366 -230 -332
rect -2490 -393 -760 -390
rect -2974 -434 -2940 -400
rect -2906 -434 -2873 -400
rect -2974 -468 -2873 -434
rect -2974 -502 -2940 -468
rect -2906 -502 -2873 -468
rect -2974 -702 -2873 -502
rect -2974 -736 -2940 -702
rect -2906 -736 -2873 -702
rect -2974 -770 -2873 -736
rect -2974 -804 -2940 -770
rect -2906 -804 -2873 -770
rect -2974 -838 -2873 -804
rect -2811 -400 -393 -393
rect -2811 -417 -2298 -400
rect -2811 -451 -2787 -417
rect -2753 -451 -2719 -417
rect -2685 -451 -2519 -417
rect -2485 -451 -2451 -417
rect -2417 -434 -2298 -417
rect -2264 -434 -1940 -400
rect -1906 -417 -1298 -400
rect -1906 -434 -1787 -417
rect -2417 -451 -1787 -434
rect -1753 -451 -1719 -417
rect -1685 -451 -1519 -417
rect -1485 -451 -1451 -417
rect -1417 -434 -1298 -417
rect -1264 -434 -940 -400
rect -906 -417 -393 -400
rect -906 -434 -787 -417
rect -1417 -451 -787 -434
rect -753 -451 -719 -417
rect -685 -451 -519 -417
rect -485 -451 -451 -417
rect -417 -451 -393 -417
rect -2811 -460 -393 -451
rect -2811 -465 -2393 -460
rect -2811 -485 -2739 -465
rect -2811 -519 -2787 -485
rect -2753 -519 -2739 -485
rect -2811 -685 -2739 -519
rect -2465 -485 -2393 -465
rect -2465 -519 -2451 -485
rect -2417 -519 -2393 -485
rect -2681 -537 -2523 -523
rect -2681 -571 -2667 -537
rect -2633 -551 -2571 -537
rect -2537 -571 -2523 -537
rect -2681 -633 -2653 -571
rect -2551 -633 -2523 -571
rect -2681 -667 -2667 -633
rect -2633 -667 -2571 -653
rect -2537 -667 -2523 -633
rect -2681 -681 -2523 -667
rect -2811 -719 -2787 -685
rect -2753 -719 -2739 -685
rect -2811 -739 -2739 -719
rect -2465 -685 -2393 -519
rect -2465 -719 -2451 -685
rect -2417 -719 -2393 -685
rect -2465 -739 -2393 -719
rect -2811 -753 -2393 -739
rect -2811 -787 -2787 -753
rect -2753 -787 -2719 -753
rect -2685 -787 -2519 -753
rect -2485 -787 -2451 -753
rect -2417 -787 -2393 -753
rect -2811 -811 -2393 -787
rect -2331 -468 -2230 -460
rect -2331 -502 -2298 -468
rect -2264 -502 -2230 -468
rect -2331 -702 -2230 -502
rect -2331 -736 -2298 -702
rect -2264 -736 -2230 -702
rect -2331 -770 -2230 -736
rect -2331 -804 -2298 -770
rect -2264 -804 -2230 -770
rect -2974 -872 -2940 -838
rect -2906 -872 -2873 -838
rect -2974 -873 -2873 -872
rect -2331 -838 -2230 -804
rect -2331 -872 -2298 -838
rect -2264 -872 -2230 -838
rect -2331 -873 -2230 -872
rect -2974 -906 -2230 -873
rect -2974 -940 -2940 -906
rect -2906 -940 -2872 -906
rect -2838 -940 -2804 -906
rect -2770 -940 -2736 -906
rect -2702 -940 -2502 -906
rect -2468 -940 -2434 -906
rect -2400 -940 -2366 -906
rect -2332 -940 -2298 -906
rect -2264 -940 -2230 -906
rect -2974 -974 -2230 -940
rect -2120 -1230 -2080 -460
rect -1974 -468 -1873 -460
rect -1974 -502 -1940 -468
rect -1906 -502 -1873 -468
rect -1974 -702 -1873 -502
rect -1974 -736 -1940 -702
rect -1906 -736 -1873 -702
rect -1974 -770 -1873 -736
rect -1974 -804 -1940 -770
rect -1906 -804 -1873 -770
rect -1974 -838 -1873 -804
rect -1811 -465 -1393 -460
rect -1811 -485 -1739 -465
rect -1811 -519 -1787 -485
rect -1753 -519 -1739 -485
rect -1811 -685 -1739 -519
rect -1465 -485 -1393 -465
rect -1465 -519 -1451 -485
rect -1417 -519 -1393 -485
rect -1681 -537 -1523 -523
rect -1681 -571 -1667 -537
rect -1633 -551 -1571 -537
rect -1537 -571 -1523 -537
rect -1681 -633 -1653 -571
rect -1551 -633 -1523 -571
rect -1681 -667 -1667 -633
rect -1633 -667 -1571 -653
rect -1537 -667 -1523 -633
rect -1681 -681 -1523 -667
rect -1811 -719 -1787 -685
rect -1753 -719 -1739 -685
rect -1811 -739 -1739 -719
rect -1465 -685 -1393 -519
rect -1465 -719 -1451 -685
rect -1417 -719 -1393 -685
rect -1465 -739 -1393 -719
rect -1811 -753 -1393 -739
rect -1811 -787 -1787 -753
rect -1753 -787 -1719 -753
rect -1685 -787 -1519 -753
rect -1485 -787 -1451 -753
rect -1417 -787 -1393 -753
rect -1811 -811 -1393 -787
rect -1331 -468 -1230 -460
rect -1331 -502 -1298 -468
rect -1264 -502 -1230 -468
rect -1331 -702 -1230 -502
rect -1331 -736 -1298 -702
rect -1264 -736 -1230 -702
rect -1331 -770 -1230 -736
rect -1331 -804 -1298 -770
rect -1264 -804 -1230 -770
rect -1974 -872 -1940 -838
rect -1906 -872 -1873 -838
rect -1974 -873 -1873 -872
rect -1331 -838 -1230 -804
rect -1331 -872 -1298 -838
rect -1264 -872 -1230 -838
rect -1331 -873 -1230 -872
rect -1974 -880 -1230 -873
rect -974 -468 -873 -460
rect -974 -502 -940 -468
rect -906 -502 -873 -468
rect -974 -702 -873 -502
rect -974 -736 -940 -702
rect -906 -736 -873 -702
rect -974 -770 -873 -736
rect -974 -804 -940 -770
rect -906 -804 -873 -770
rect -974 -838 -873 -804
rect -811 -465 -393 -460
rect -811 -485 -739 -465
rect -811 -519 -787 -485
rect -753 -519 -739 -485
rect -811 -685 -739 -519
rect -465 -485 -393 -465
rect -465 -519 -451 -485
rect -417 -519 -393 -485
rect -681 -537 -523 -523
rect -681 -571 -667 -537
rect -633 -551 -571 -537
rect -537 -571 -523 -537
rect -681 -633 -653 -571
rect -551 -633 -523 -571
rect -681 -667 -667 -633
rect -633 -667 -571 -653
rect -537 -667 -523 -633
rect -681 -681 -523 -667
rect -811 -719 -787 -685
rect -753 -719 -739 -685
rect -811 -739 -739 -719
rect -465 -685 -393 -519
rect -465 -719 -451 -685
rect -417 -719 -393 -685
rect -465 -739 -393 -719
rect -811 -753 -393 -739
rect -811 -787 -787 -753
rect -753 -787 -719 -753
rect -685 -787 -519 -753
rect -485 -787 -451 -753
rect -417 -787 -393 -753
rect -811 -811 -393 -787
rect -331 -400 -230 -366
rect -331 -434 -298 -400
rect -264 -434 -230 -400
rect -331 -468 -230 -434
rect -331 -502 -298 -468
rect -264 -502 -230 -468
rect -331 -702 -230 -502
rect -331 -736 -298 -702
rect -264 -736 -230 -702
rect -331 -770 -230 -736
rect -331 -804 -298 -770
rect -264 -804 -230 -770
rect -974 -872 -940 -838
rect -906 -872 -873 -838
rect -974 -873 -873 -872
rect -331 -838 -230 -804
rect -331 -872 -298 -838
rect -264 -872 -230 -838
rect -331 -873 -230 -872
rect -974 -880 -230 -873
rect -1974 -906 -230 -880
rect -1974 -940 -1940 -906
rect -1906 -940 -1872 -906
rect -1838 -940 -1804 -906
rect -1770 -940 -1736 -906
rect -1702 -940 -1502 -906
rect -1468 -940 -1434 -906
rect -1400 -940 -1366 -906
rect -1332 -940 -1298 -906
rect -1264 -940 -940 -906
rect -906 -940 -872 -906
rect -838 -940 -804 -906
rect -770 -940 -736 -906
rect -702 -940 -502 -906
rect -468 -940 -434 -906
rect -400 -940 -366 -906
rect -332 -940 -298 -906
rect -264 -940 -230 -906
rect -1974 -970 -230 -940
rect -1974 -974 -1230 -970
rect -974 -974 -230 -970
rect 26 -264 770 -230
rect 26 -298 60 -264
rect 94 -298 128 -264
rect 162 -298 196 -264
rect 230 -298 264 -264
rect 298 -298 498 -264
rect 532 -298 566 -264
rect 600 -298 634 -264
rect 668 -298 702 -264
rect 736 -298 770 -264
rect 26 -331 770 -298
rect 26 -332 127 -331
rect 26 -366 60 -332
rect 94 -366 127 -332
rect 26 -400 127 -366
rect 669 -332 770 -331
rect 669 -366 702 -332
rect 736 -366 770 -332
rect 26 -434 60 -400
rect 94 -434 127 -400
rect 26 -468 127 -434
rect 26 -502 60 -468
rect 94 -502 127 -468
rect 26 -702 127 -502
rect 26 -736 60 -702
rect 94 -736 127 -702
rect 26 -770 127 -736
rect 26 -804 60 -770
rect 94 -804 127 -770
rect 26 -838 127 -804
rect 189 -417 607 -393
rect 189 -451 213 -417
rect 247 -451 281 -417
rect 315 -451 481 -417
rect 515 -451 549 -417
rect 583 -451 607 -417
rect 189 -465 607 -451
rect 189 -485 261 -465
rect 189 -519 213 -485
rect 247 -519 261 -485
rect 189 -685 261 -519
rect 535 -485 607 -465
rect 535 -519 549 -485
rect 583 -519 607 -485
rect 319 -537 477 -523
rect 319 -571 333 -537
rect 367 -551 429 -537
rect 463 -571 477 -537
rect 319 -633 347 -571
rect 449 -633 477 -571
rect 319 -667 333 -633
rect 367 -667 429 -653
rect 463 -667 477 -633
rect 319 -681 477 -667
rect 189 -719 213 -685
rect 247 -719 261 -685
rect 189 -739 261 -719
rect 535 -685 607 -519
rect 535 -719 549 -685
rect 583 -719 607 -685
rect 535 -739 607 -719
rect 189 -753 607 -739
rect 189 -787 213 -753
rect 247 -787 281 -753
rect 315 -787 481 -753
rect 515 -787 549 -753
rect 583 -787 607 -753
rect 189 -811 607 -787
rect 669 -400 770 -366
rect 669 -434 702 -400
rect 736 -434 770 -400
rect 669 -468 770 -434
rect 669 -502 702 -468
rect 736 -502 770 -468
rect 669 -702 770 -502
rect 669 -736 702 -702
rect 736 -736 770 -702
rect 669 -770 770 -736
rect 669 -804 702 -770
rect 736 -804 770 -770
rect 26 -872 60 -838
rect 94 -872 127 -838
rect 26 -873 127 -872
rect 190 -873 260 -811
rect 669 -838 770 -804
rect 669 -872 702 -838
rect 736 -872 770 -838
rect 669 -873 770 -872
rect 26 -906 770 -873
rect 26 -940 60 -906
rect 94 -940 128 -906
rect 162 -940 196 -906
rect 230 -940 264 -906
rect 298 -940 498 -906
rect 532 -940 566 -906
rect 600 -940 634 -906
rect 668 -940 702 -906
rect 736 -940 770 -906
rect 26 -974 770 -940
rect 1026 -264 1770 -230
rect 1026 -298 1060 -264
rect 1094 -298 1128 -264
rect 1162 -298 1196 -264
rect 1230 -298 1264 -264
rect 1298 -298 1498 -264
rect 1532 -298 1566 -264
rect 1600 -298 1634 -264
rect 1668 -298 1702 -264
rect 1736 -298 1770 -264
rect 1026 -331 1770 -298
rect 1026 -332 1127 -331
rect 1026 -366 1060 -332
rect 1094 -366 1127 -332
rect 1026 -400 1127 -366
rect 1669 -332 1770 -331
rect 1669 -366 1702 -332
rect 1736 -366 1770 -332
rect 1026 -434 1060 -400
rect 1094 -434 1127 -400
rect 1026 -468 1127 -434
rect 1026 -502 1060 -468
rect 1094 -502 1127 -468
rect 1026 -702 1127 -502
rect 1026 -736 1060 -702
rect 1094 -736 1127 -702
rect 1026 -770 1127 -736
rect 1026 -804 1060 -770
rect 1094 -804 1127 -770
rect 1026 -838 1127 -804
rect 1189 -417 1607 -393
rect 1189 -451 1213 -417
rect 1247 -451 1281 -417
rect 1315 -451 1481 -417
rect 1515 -451 1549 -417
rect 1583 -451 1607 -417
rect 1189 -465 1607 -451
rect 1189 -485 1261 -465
rect 1189 -519 1213 -485
rect 1247 -519 1261 -485
rect 1189 -685 1261 -519
rect 1535 -485 1607 -465
rect 1535 -519 1549 -485
rect 1583 -519 1607 -485
rect 1319 -537 1477 -523
rect 1319 -571 1333 -537
rect 1367 -551 1429 -537
rect 1463 -571 1477 -537
rect 1319 -633 1347 -571
rect 1449 -633 1477 -571
rect 1319 -667 1333 -633
rect 1367 -667 1429 -653
rect 1463 -667 1477 -633
rect 1319 -681 1477 -667
rect 1189 -719 1213 -685
rect 1247 -719 1261 -685
rect 1189 -739 1261 -719
rect 1535 -685 1607 -519
rect 1535 -719 1549 -685
rect 1583 -719 1607 -685
rect 1535 -739 1607 -719
rect 1189 -753 1607 -739
rect 1189 -787 1213 -753
rect 1247 -787 1281 -753
rect 1315 -787 1481 -753
rect 1515 -787 1549 -753
rect 1583 -787 1607 -753
rect 1189 -811 1607 -787
rect 1669 -400 1770 -366
rect 1669 -434 1702 -400
rect 1736 -434 1770 -400
rect 1669 -468 1770 -434
rect 1669 -502 1702 -468
rect 1736 -502 1770 -468
rect 1669 -702 1770 -502
rect 1669 -736 1702 -702
rect 1736 -736 1770 -702
rect 1669 -770 1770 -736
rect 1669 -804 1702 -770
rect 1736 -804 1770 -770
rect 1026 -872 1060 -838
rect 1094 -872 1127 -838
rect 1026 -873 1127 -872
rect 1669 -838 1770 -804
rect 1669 -872 1702 -838
rect 1736 -872 1770 -838
rect 1669 -873 1770 -872
rect 1026 -906 1770 -873
rect 1026 -940 1060 -906
rect 1094 -940 1128 -906
rect 1162 -940 1196 -906
rect 1230 -940 1264 -906
rect 1298 -940 1498 -906
rect 1532 -940 1566 -906
rect 1600 -940 1634 -906
rect 1668 -940 1702 -906
rect 1736 -940 1770 -906
rect 1026 -974 1770 -940
rect -1330 -1230 -1230 -974
rect -3974 -1264 -3230 -1230
rect -3974 -1298 -3940 -1264
rect -3906 -1298 -3872 -1264
rect -3838 -1298 -3804 -1264
rect -3770 -1298 -3736 -1264
rect -3702 -1298 -3502 -1264
rect -3468 -1298 -3434 -1264
rect -3400 -1298 -3366 -1264
rect -3332 -1298 -3298 -1264
rect -3264 -1298 -3230 -1264
rect -3974 -1331 -3230 -1298
rect -3974 -1332 -3873 -1331
rect -3974 -1366 -3940 -1332
rect -3906 -1366 -3873 -1332
rect -3974 -1400 -3873 -1366
rect -3331 -1332 -3230 -1331
rect -3331 -1366 -3298 -1332
rect -3264 -1366 -3230 -1332
rect -3974 -1434 -3940 -1400
rect -3906 -1434 -3873 -1400
rect -3974 -1468 -3873 -1434
rect -3974 -1502 -3940 -1468
rect -3906 -1502 -3873 -1468
rect -3974 -1702 -3873 -1502
rect -3974 -1736 -3940 -1702
rect -3906 -1736 -3873 -1702
rect -3974 -1770 -3873 -1736
rect -3974 -1804 -3940 -1770
rect -3906 -1804 -3873 -1770
rect -3974 -1838 -3873 -1804
rect -3811 -1417 -3393 -1393
rect -3811 -1451 -3787 -1417
rect -3753 -1451 -3719 -1417
rect -3685 -1451 -3519 -1417
rect -3485 -1451 -3451 -1417
rect -3417 -1451 -3393 -1417
rect -3811 -1465 -3393 -1451
rect -3811 -1485 -3739 -1465
rect -3811 -1519 -3787 -1485
rect -3753 -1519 -3739 -1485
rect -3811 -1685 -3739 -1519
rect -3465 -1485 -3393 -1465
rect -3465 -1519 -3451 -1485
rect -3417 -1519 -3393 -1485
rect -3681 -1537 -3523 -1523
rect -3681 -1571 -3667 -1537
rect -3633 -1551 -3571 -1537
rect -3537 -1571 -3523 -1537
rect -3681 -1633 -3653 -1571
rect -3551 -1633 -3523 -1571
rect -3681 -1667 -3667 -1633
rect -3633 -1667 -3571 -1653
rect -3537 -1667 -3523 -1633
rect -3681 -1681 -3523 -1667
rect -3811 -1719 -3787 -1685
rect -3753 -1719 -3739 -1685
rect -3811 -1739 -3739 -1719
rect -3465 -1685 -3393 -1519
rect -3465 -1719 -3451 -1685
rect -3417 -1719 -3393 -1685
rect -3465 -1739 -3393 -1719
rect -3811 -1753 -3393 -1739
rect -3811 -1787 -3787 -1753
rect -3753 -1787 -3719 -1753
rect -3685 -1787 -3519 -1753
rect -3485 -1787 -3451 -1753
rect -3417 -1787 -3393 -1753
rect -3811 -1811 -3393 -1787
rect -3331 -1400 -3230 -1366
rect -3331 -1434 -3298 -1400
rect -3264 -1434 -3230 -1400
rect -3331 -1468 -3230 -1434
rect -3331 -1502 -3298 -1468
rect -3264 -1502 -3230 -1468
rect -3331 -1702 -3230 -1502
rect -3331 -1736 -3298 -1702
rect -3264 -1736 -3230 -1702
rect -3331 -1770 -3230 -1736
rect -3331 -1804 -3298 -1770
rect -3264 -1804 -3230 -1770
rect -3974 -1872 -3940 -1838
rect -3906 -1872 -3873 -1838
rect -3974 -1873 -3873 -1872
rect -3331 -1838 -3230 -1804
rect -3331 -1872 -3298 -1838
rect -3264 -1872 -3230 -1838
rect -3331 -1873 -3230 -1872
rect -3974 -1906 -3230 -1873
rect -3974 -1940 -3940 -1906
rect -3906 -1940 -3872 -1906
rect -3838 -1940 -3804 -1906
rect -3770 -1940 -3736 -1906
rect -3702 -1940 -3502 -1906
rect -3468 -1940 -3434 -1906
rect -3400 -1940 -3366 -1906
rect -3332 -1940 -3298 -1906
rect -3264 -1940 -3230 -1906
rect -3974 -1974 -3230 -1940
rect -2974 -1264 -1230 -1230
rect -2974 -1298 -2940 -1264
rect -2906 -1298 -2872 -1264
rect -2838 -1298 -2804 -1264
rect -2770 -1298 -2736 -1264
rect -2702 -1298 -2502 -1264
rect -2468 -1298 -2434 -1264
rect -2400 -1298 -2366 -1264
rect -2332 -1298 -2298 -1264
rect -2264 -1298 -1940 -1264
rect -1906 -1298 -1872 -1264
rect -1838 -1298 -1804 -1264
rect -1770 -1298 -1736 -1264
rect -1702 -1298 -1502 -1264
rect -1468 -1298 -1434 -1264
rect -1400 -1298 -1366 -1264
rect -1332 -1298 -1298 -1264
rect -1264 -1298 -1230 -1264
rect -2974 -1330 -1230 -1298
rect -2974 -1331 -2230 -1330
rect -2974 -1332 -2873 -1331
rect -2974 -1366 -2940 -1332
rect -2906 -1366 -2873 -1332
rect -2974 -1400 -2873 -1366
rect -2331 -1332 -2230 -1331
rect -2331 -1366 -2298 -1332
rect -2264 -1366 -2230 -1332
rect -2331 -1390 -2230 -1366
rect -2120 -1390 -2080 -1330
rect -1974 -1331 -1230 -1330
rect -1974 -1332 -1873 -1331
rect -1974 -1366 -1940 -1332
rect -1906 -1366 -1873 -1332
rect -1974 -1390 -1873 -1366
rect -1331 -1332 -1230 -1331
rect -1331 -1366 -1298 -1332
rect -1264 -1366 -1230 -1332
rect -2480 -1393 -1790 -1390
rect -2974 -1434 -2940 -1400
rect -2906 -1434 -2873 -1400
rect -2974 -1468 -2873 -1434
rect -2974 -1502 -2940 -1468
rect -2906 -1502 -2873 -1468
rect -2974 -1702 -2873 -1502
rect -2974 -1736 -2940 -1702
rect -2906 -1736 -2873 -1702
rect -2974 -1770 -2873 -1736
rect -2974 -1804 -2940 -1770
rect -2906 -1804 -2873 -1770
rect -2974 -1838 -2873 -1804
rect -2811 -1400 -1393 -1393
rect -2811 -1417 -2298 -1400
rect -2811 -1451 -2787 -1417
rect -2753 -1451 -2719 -1417
rect -2685 -1451 -2519 -1417
rect -2485 -1451 -2451 -1417
rect -2417 -1434 -2298 -1417
rect -2264 -1434 -1940 -1400
rect -1906 -1417 -1393 -1400
rect -1906 -1434 -1787 -1417
rect -2417 -1451 -1787 -1434
rect -1753 -1451 -1719 -1417
rect -1685 -1451 -1519 -1417
rect -1485 -1451 -1451 -1417
rect -1417 -1451 -1393 -1417
rect -2811 -1465 -1393 -1451
rect -2811 -1485 -2739 -1465
rect -2480 -1468 -1739 -1465
rect -2480 -1470 -2298 -1468
rect -2811 -1519 -2787 -1485
rect -2753 -1519 -2739 -1485
rect -2811 -1685 -2739 -1519
rect -2465 -1485 -2393 -1470
rect -2465 -1519 -2451 -1485
rect -2417 -1519 -2393 -1485
rect -2681 -1537 -2523 -1523
rect -2681 -1571 -2667 -1537
rect -2633 -1551 -2571 -1537
rect -2537 -1571 -2523 -1537
rect -2681 -1633 -2653 -1571
rect -2551 -1633 -2523 -1571
rect -2681 -1667 -2667 -1633
rect -2633 -1667 -2571 -1653
rect -2537 -1667 -2523 -1633
rect -2681 -1681 -2523 -1667
rect -2811 -1719 -2787 -1685
rect -2753 -1719 -2739 -1685
rect -2811 -1739 -2739 -1719
rect -2465 -1685 -2393 -1519
rect -2465 -1719 -2451 -1685
rect -2417 -1719 -2393 -1685
rect -2465 -1739 -2393 -1719
rect -2811 -1753 -2393 -1739
rect -2811 -1787 -2787 -1753
rect -2753 -1787 -2719 -1753
rect -2685 -1787 -2519 -1753
rect -2485 -1787 -2451 -1753
rect -2417 -1787 -2393 -1753
rect -2811 -1811 -2393 -1787
rect -2331 -1502 -2298 -1470
rect -2264 -1470 -1940 -1468
rect -2264 -1502 -2230 -1470
rect -2331 -1702 -2230 -1502
rect -2331 -1736 -2298 -1702
rect -2264 -1736 -2230 -1702
rect -2331 -1770 -2230 -1736
rect -2331 -1804 -2298 -1770
rect -2264 -1804 -2230 -1770
rect -2974 -1872 -2940 -1838
rect -2906 -1872 -2873 -1838
rect -2974 -1873 -2873 -1872
rect -2331 -1838 -2230 -1804
rect -2331 -1872 -2298 -1838
rect -2264 -1872 -2230 -1838
rect -2331 -1873 -2230 -1872
rect -2974 -1906 -2230 -1873
rect -2974 -1940 -2940 -1906
rect -2906 -1940 -2872 -1906
rect -2838 -1940 -2804 -1906
rect -2770 -1940 -2736 -1906
rect -2702 -1940 -2502 -1906
rect -2468 -1940 -2434 -1906
rect -2400 -1940 -2366 -1906
rect -2332 -1940 -2298 -1906
rect -2264 -1940 -2230 -1906
rect -2974 -1974 -2230 -1940
rect -1974 -1502 -1940 -1470
rect -1906 -1470 -1739 -1468
rect -1906 -1502 -1873 -1470
rect -1974 -1702 -1873 -1502
rect -1974 -1736 -1940 -1702
rect -1906 -1736 -1873 -1702
rect -1974 -1770 -1873 -1736
rect -1974 -1804 -1940 -1770
rect -1906 -1804 -1873 -1770
rect -1974 -1838 -1873 -1804
rect -1811 -1485 -1739 -1470
rect -1811 -1519 -1787 -1485
rect -1753 -1519 -1739 -1485
rect -1811 -1685 -1739 -1519
rect -1465 -1485 -1393 -1465
rect -1465 -1519 -1451 -1485
rect -1417 -1519 -1393 -1485
rect -1681 -1537 -1523 -1523
rect -1681 -1571 -1667 -1537
rect -1633 -1551 -1571 -1537
rect -1537 -1571 -1523 -1537
rect -1681 -1633 -1653 -1571
rect -1551 -1633 -1523 -1571
rect -1681 -1667 -1667 -1633
rect -1633 -1667 -1571 -1653
rect -1537 -1667 -1523 -1633
rect -1681 -1681 -1523 -1667
rect -1811 -1719 -1787 -1685
rect -1753 -1719 -1739 -1685
rect -1811 -1739 -1739 -1719
rect -1465 -1685 -1393 -1519
rect -1465 -1719 -1451 -1685
rect -1417 -1719 -1393 -1685
rect -1465 -1739 -1393 -1719
rect -1811 -1753 -1393 -1739
rect -1811 -1787 -1787 -1753
rect -1753 -1787 -1719 -1753
rect -1685 -1787 -1519 -1753
rect -1485 -1787 -1451 -1753
rect -1417 -1787 -1393 -1753
rect -1811 -1811 -1393 -1787
rect -1331 -1400 -1230 -1366
rect -1331 -1434 -1298 -1400
rect -1264 -1434 -1230 -1400
rect -1331 -1468 -1230 -1434
rect -1331 -1502 -1298 -1468
rect -1264 -1502 -1230 -1468
rect -1331 -1702 -1230 -1502
rect -1331 -1736 -1298 -1702
rect -1264 -1736 -1230 -1702
rect -1331 -1770 -1230 -1736
rect -1331 -1804 -1298 -1770
rect -1264 -1804 -1230 -1770
rect -1974 -1872 -1940 -1838
rect -1906 -1872 -1873 -1838
rect -1974 -1873 -1873 -1872
rect -1331 -1838 -1230 -1804
rect -1331 -1872 -1298 -1838
rect -1264 -1872 -1230 -1838
rect -1331 -1873 -1230 -1872
rect -1974 -1906 -1230 -1873
rect -1974 -1940 -1940 -1906
rect -1906 -1940 -1872 -1906
rect -1838 -1940 -1804 -1906
rect -1770 -1940 -1736 -1906
rect -1702 -1940 -1502 -1906
rect -1468 -1940 -1434 -1906
rect -1400 -1940 -1366 -1906
rect -1332 -1940 -1298 -1906
rect -1264 -1940 -1230 -1906
rect -1974 -1974 -1230 -1940
rect -974 -1264 -230 -1230
rect -974 -1298 -940 -1264
rect -906 -1298 -872 -1264
rect -838 -1298 -804 -1264
rect -770 -1298 -736 -1264
rect -702 -1298 -502 -1264
rect -468 -1298 -434 -1264
rect -400 -1298 -366 -1264
rect -332 -1298 -298 -1264
rect -264 -1298 -230 -1264
rect -974 -1331 -230 -1298
rect -974 -1332 -873 -1331
rect -974 -1366 -940 -1332
rect -906 -1366 -873 -1332
rect -974 -1400 -873 -1366
rect -331 -1332 -230 -1331
rect -331 -1366 -298 -1332
rect -264 -1366 -230 -1332
rect -974 -1434 -940 -1400
rect -906 -1434 -873 -1400
rect -974 -1468 -873 -1434
rect -974 -1502 -940 -1468
rect -906 -1502 -873 -1468
rect -974 -1702 -873 -1502
rect -974 -1736 -940 -1702
rect -906 -1736 -873 -1702
rect -974 -1770 -873 -1736
rect -974 -1804 -940 -1770
rect -906 -1804 -873 -1770
rect -974 -1838 -873 -1804
rect -811 -1417 -393 -1393
rect -811 -1451 -787 -1417
rect -753 -1451 -719 -1417
rect -685 -1451 -519 -1417
rect -485 -1451 -451 -1417
rect -417 -1451 -393 -1417
rect -811 -1465 -393 -1451
rect -811 -1485 -739 -1465
rect -811 -1519 -787 -1485
rect -753 -1519 -739 -1485
rect -811 -1685 -739 -1519
rect -465 -1485 -393 -1465
rect -465 -1519 -451 -1485
rect -417 -1519 -393 -1485
rect -681 -1537 -523 -1523
rect -681 -1571 -667 -1537
rect -633 -1551 -571 -1537
rect -537 -1571 -523 -1537
rect -681 -1633 -653 -1571
rect -551 -1633 -523 -1571
rect -681 -1667 -667 -1633
rect -633 -1667 -571 -1653
rect -537 -1667 -523 -1633
rect -681 -1681 -523 -1667
rect -811 -1719 -787 -1685
rect -753 -1719 -739 -1685
rect -811 -1739 -739 -1719
rect -465 -1685 -393 -1519
rect -465 -1719 -451 -1685
rect -417 -1719 -393 -1685
rect -465 -1739 -393 -1719
rect -811 -1753 -393 -1739
rect -811 -1787 -787 -1753
rect -753 -1787 -719 -1753
rect -685 -1787 -519 -1753
rect -485 -1787 -451 -1753
rect -417 -1787 -393 -1753
rect -811 -1811 -393 -1787
rect -331 -1400 -230 -1366
rect -331 -1434 -298 -1400
rect -264 -1434 -230 -1400
rect -331 -1468 -230 -1434
rect -331 -1502 -298 -1468
rect -264 -1502 -230 -1468
rect -331 -1702 -230 -1502
rect -331 -1736 -298 -1702
rect -264 -1736 -230 -1702
rect -331 -1770 -230 -1736
rect -331 -1804 -298 -1770
rect -264 -1804 -230 -1770
rect -974 -1872 -940 -1838
rect -906 -1872 -873 -1838
rect -974 -1873 -873 -1872
rect -810 -1873 -740 -1811
rect -331 -1838 -230 -1804
rect -331 -1872 -298 -1838
rect -264 -1872 -230 -1838
rect -331 -1873 -230 -1872
rect -974 -1906 -230 -1873
rect -974 -1940 -940 -1906
rect -906 -1940 -872 -1906
rect -838 -1940 -804 -1906
rect -770 -1940 -736 -1906
rect -702 -1940 -502 -1906
rect -468 -1940 -434 -1906
rect -400 -1940 -366 -1906
rect -332 -1940 -298 -1906
rect -264 -1940 -230 -1906
rect -974 -1974 -230 -1940
rect 26 -1264 770 -1230
rect 26 -1298 60 -1264
rect 94 -1298 128 -1264
rect 162 -1298 196 -1264
rect 230 -1298 264 -1264
rect 298 -1298 498 -1264
rect 532 -1298 566 -1264
rect 600 -1298 634 -1264
rect 668 -1298 702 -1264
rect 736 -1298 770 -1264
rect 26 -1331 770 -1298
rect 26 -1332 127 -1331
rect 26 -1366 60 -1332
rect 94 -1366 127 -1332
rect 26 -1400 127 -1366
rect 669 -1332 770 -1331
rect 669 -1366 702 -1332
rect 736 -1366 770 -1332
rect 26 -1434 60 -1400
rect 94 -1434 127 -1400
rect 26 -1468 127 -1434
rect 26 -1502 60 -1468
rect 94 -1502 127 -1468
rect 26 -1702 127 -1502
rect 26 -1736 60 -1702
rect 94 -1736 127 -1702
rect 26 -1770 127 -1736
rect 26 -1804 60 -1770
rect 94 -1804 127 -1770
rect 26 -1838 127 -1804
rect 189 -1410 607 -1393
rect 189 -1417 550 -1410
rect 189 -1451 213 -1417
rect 247 -1451 281 -1417
rect 315 -1451 481 -1417
rect 515 -1451 549 -1417
rect 590 -1450 607 -1410
rect 583 -1451 607 -1450
rect 189 -1465 607 -1451
rect 189 -1485 261 -1465
rect 189 -1519 213 -1485
rect 247 -1519 261 -1485
rect 189 -1685 261 -1519
rect 535 -1485 607 -1465
rect 535 -1519 549 -1485
rect 583 -1519 607 -1485
rect 319 -1537 477 -1523
rect 319 -1571 333 -1537
rect 367 -1551 429 -1537
rect 463 -1571 477 -1537
rect 319 -1633 347 -1571
rect 449 -1633 477 -1571
rect 319 -1667 333 -1633
rect 367 -1667 429 -1653
rect 463 -1667 477 -1633
rect 319 -1681 477 -1667
rect 189 -1719 213 -1685
rect 247 -1719 261 -1685
rect 189 -1739 261 -1719
rect 535 -1685 607 -1519
rect 535 -1719 549 -1685
rect 583 -1719 607 -1685
rect 535 -1739 607 -1719
rect 189 -1753 607 -1739
rect 189 -1787 213 -1753
rect 247 -1787 281 -1753
rect 315 -1787 481 -1753
rect 515 -1787 549 -1753
rect 583 -1787 607 -1753
rect 189 -1811 607 -1787
rect 669 -1400 770 -1366
rect 669 -1434 702 -1400
rect 736 -1434 770 -1400
rect 669 -1468 770 -1434
rect 669 -1502 702 -1468
rect 736 -1502 770 -1468
rect 669 -1702 770 -1502
rect 669 -1736 702 -1702
rect 736 -1736 770 -1702
rect 669 -1770 770 -1736
rect 669 -1804 702 -1770
rect 736 -1804 770 -1770
rect 26 -1872 60 -1838
rect 94 -1872 127 -1838
rect 26 -1873 127 -1872
rect 669 -1838 770 -1804
rect 669 -1872 702 -1838
rect 736 -1872 770 -1838
rect 669 -1873 770 -1872
rect 26 -1900 770 -1873
rect 26 -1906 700 -1900
rect 26 -1940 60 -1906
rect 94 -1940 128 -1906
rect 162 -1940 196 -1906
rect 230 -1940 264 -1906
rect 298 -1940 498 -1906
rect 532 -1940 566 -1906
rect 600 -1940 634 -1906
rect 668 -1940 700 -1906
rect 740 -1940 770 -1900
rect 26 -1974 770 -1940
rect 1026 -1264 1770 -1230
rect 1026 -1298 1060 -1264
rect 1094 -1298 1128 -1264
rect 1162 -1298 1196 -1264
rect 1230 -1298 1264 -1264
rect 1298 -1298 1498 -1264
rect 1532 -1298 1566 -1264
rect 1600 -1298 1634 -1264
rect 1668 -1298 1702 -1264
rect 1736 -1298 1770 -1264
rect 1026 -1331 1770 -1298
rect 1026 -1332 1127 -1331
rect 1026 -1366 1060 -1332
rect 1094 -1366 1127 -1332
rect 1026 -1400 1127 -1366
rect 1669 -1332 1770 -1331
rect 1669 -1366 1702 -1332
rect 1736 -1366 1770 -1332
rect 1026 -1434 1060 -1400
rect 1094 -1434 1127 -1400
rect 1026 -1468 1127 -1434
rect 1026 -1502 1060 -1468
rect 1094 -1502 1127 -1468
rect 1026 -1702 1127 -1502
rect 1026 -1736 1060 -1702
rect 1094 -1736 1127 -1702
rect 1026 -1770 1127 -1736
rect 1026 -1804 1060 -1770
rect 1094 -1804 1127 -1770
rect 1026 -1838 1127 -1804
rect 1189 -1417 1607 -1393
rect 1189 -1451 1213 -1417
rect 1247 -1451 1281 -1417
rect 1315 -1451 1481 -1417
rect 1515 -1451 1549 -1417
rect 1583 -1451 1607 -1417
rect 1189 -1465 1607 -1451
rect 1189 -1485 1261 -1465
rect 1189 -1519 1213 -1485
rect 1247 -1519 1261 -1485
rect 1189 -1685 1261 -1519
rect 1535 -1485 1607 -1465
rect 1535 -1519 1549 -1485
rect 1583 -1519 1607 -1485
rect 1319 -1537 1477 -1523
rect 1319 -1571 1333 -1537
rect 1367 -1551 1429 -1537
rect 1463 -1571 1477 -1537
rect 1319 -1633 1347 -1571
rect 1449 -1633 1477 -1571
rect 1319 -1667 1333 -1633
rect 1367 -1667 1429 -1653
rect 1463 -1667 1477 -1633
rect 1319 -1681 1477 -1667
rect 1189 -1719 1213 -1685
rect 1247 -1719 1261 -1685
rect 1189 -1739 1261 -1719
rect 1535 -1685 1607 -1519
rect 1535 -1719 1549 -1685
rect 1583 -1719 1607 -1685
rect 1535 -1739 1607 -1719
rect 1189 -1753 1607 -1739
rect 1189 -1787 1213 -1753
rect 1247 -1787 1281 -1753
rect 1315 -1787 1481 -1753
rect 1515 -1787 1549 -1753
rect 1583 -1787 1607 -1753
rect 1189 -1811 1607 -1787
rect 1669 -1400 1770 -1366
rect 1669 -1434 1702 -1400
rect 1736 -1434 1770 -1400
rect 1669 -1468 1770 -1434
rect 1669 -1502 1702 -1468
rect 1736 -1502 1770 -1468
rect 1669 -1702 1770 -1502
rect 1669 -1736 1702 -1702
rect 1736 -1736 1770 -1702
rect 1669 -1770 1770 -1736
rect 1669 -1804 1702 -1770
rect 1736 -1804 1770 -1770
rect 1026 -1872 1060 -1838
rect 1094 -1872 1127 -1838
rect 1026 -1873 1127 -1872
rect 1669 -1838 1770 -1804
rect 1669 -1872 1702 -1838
rect 1736 -1872 1770 -1838
rect 1669 -1873 1770 -1872
rect 1026 -1906 1770 -1873
rect 1026 -1940 1060 -1906
rect 1094 -1940 1128 -1906
rect 1162 -1940 1196 -1906
rect 1230 -1940 1264 -1906
rect 1298 -1940 1498 -1906
rect 1532 -1940 1566 -1906
rect 1600 -1940 1634 -1906
rect 1668 -1940 1702 -1906
rect 1736 -1940 1770 -1906
rect 1026 -1974 1770 -1940
rect -3974 -2264 -3230 -2230
rect -3974 -2298 -3940 -2264
rect -3906 -2298 -3872 -2264
rect -3838 -2298 -3804 -2264
rect -3770 -2298 -3736 -2264
rect -3702 -2298 -3502 -2264
rect -3468 -2298 -3434 -2264
rect -3400 -2298 -3366 -2264
rect -3332 -2298 -3298 -2264
rect -3264 -2298 -3230 -2264
rect -3974 -2331 -3230 -2298
rect -3974 -2332 -3873 -2331
rect -3974 -2366 -3940 -2332
rect -3906 -2366 -3873 -2332
rect -3974 -2400 -3873 -2366
rect -3331 -2332 -3230 -2331
rect -3331 -2366 -3298 -2332
rect -3264 -2366 -3230 -2332
rect -3974 -2434 -3940 -2400
rect -3906 -2434 -3873 -2400
rect -3974 -2468 -3873 -2434
rect -3974 -2502 -3940 -2468
rect -3906 -2502 -3873 -2468
rect -3974 -2702 -3873 -2502
rect -3974 -2736 -3940 -2702
rect -3906 -2736 -3873 -2702
rect -3974 -2770 -3873 -2736
rect -3974 -2804 -3940 -2770
rect -3906 -2804 -3873 -2770
rect -3974 -2838 -3873 -2804
rect -3811 -2417 -3393 -2393
rect -3811 -2451 -3787 -2417
rect -3753 -2451 -3719 -2417
rect -3685 -2451 -3519 -2417
rect -3485 -2451 -3451 -2417
rect -3417 -2451 -3393 -2417
rect -3811 -2465 -3393 -2451
rect -3811 -2485 -3739 -2465
rect -3811 -2519 -3787 -2485
rect -3753 -2519 -3739 -2485
rect -3811 -2685 -3739 -2519
rect -3465 -2485 -3393 -2465
rect -3465 -2519 -3451 -2485
rect -3417 -2519 -3393 -2485
rect -3681 -2537 -3523 -2523
rect -3681 -2571 -3667 -2537
rect -3633 -2551 -3571 -2537
rect -3537 -2571 -3523 -2537
rect -3681 -2633 -3653 -2571
rect -3551 -2633 -3523 -2571
rect -3681 -2667 -3667 -2633
rect -3633 -2667 -3571 -2653
rect -3537 -2667 -3523 -2633
rect -3681 -2681 -3523 -2667
rect -3811 -2719 -3787 -2685
rect -3753 -2719 -3739 -2685
rect -3811 -2739 -3739 -2719
rect -3465 -2685 -3393 -2519
rect -3465 -2719 -3451 -2685
rect -3417 -2719 -3393 -2685
rect -3465 -2739 -3393 -2719
rect -3811 -2753 -3393 -2739
rect -3811 -2787 -3787 -2753
rect -3753 -2787 -3719 -2753
rect -3685 -2787 -3519 -2753
rect -3485 -2787 -3451 -2753
rect -3417 -2787 -3393 -2753
rect -3811 -2811 -3393 -2787
rect -3331 -2400 -3230 -2366
rect -3331 -2434 -3298 -2400
rect -3264 -2434 -3230 -2400
rect -3331 -2468 -3230 -2434
rect -3331 -2502 -3298 -2468
rect -3264 -2502 -3230 -2468
rect -3331 -2702 -3230 -2502
rect -3331 -2736 -3298 -2702
rect -3264 -2736 -3230 -2702
rect -3331 -2770 -3230 -2736
rect -3331 -2804 -3298 -2770
rect -3264 -2804 -3230 -2770
rect -3974 -2872 -3940 -2838
rect -3906 -2872 -3873 -2838
rect -3974 -2873 -3873 -2872
rect -3331 -2838 -3230 -2804
rect -3331 -2872 -3298 -2838
rect -3264 -2872 -3230 -2838
rect -3331 -2873 -3230 -2872
rect -3974 -2906 -3230 -2873
rect -3974 -2940 -3940 -2906
rect -3906 -2940 -3872 -2906
rect -3838 -2940 -3804 -2906
rect -3770 -2940 -3736 -2906
rect -3702 -2940 -3502 -2906
rect -3468 -2940 -3434 -2906
rect -3400 -2940 -3366 -2906
rect -3332 -2940 -3298 -2906
rect -3264 -2940 -3230 -2906
rect -3974 -2974 -3230 -2940
rect -2974 -2264 -2230 -2230
rect -2974 -2298 -2940 -2264
rect -2906 -2298 -2872 -2264
rect -2838 -2298 -2804 -2264
rect -2770 -2298 -2736 -2264
rect -2702 -2298 -2502 -2264
rect -2468 -2298 -2434 -2264
rect -2400 -2298 -2366 -2264
rect -2332 -2298 -2298 -2264
rect -2264 -2298 -2230 -2264
rect -2974 -2331 -2230 -2298
rect -2974 -2332 -2873 -2331
rect -2974 -2366 -2940 -2332
rect -2906 -2366 -2873 -2332
rect -2974 -2400 -2873 -2366
rect -2331 -2332 -2230 -2331
rect -2331 -2366 -2298 -2332
rect -2264 -2366 -2230 -2332
rect -2974 -2434 -2940 -2400
rect -2906 -2434 -2873 -2400
rect -2974 -2468 -2873 -2434
rect -2974 -2502 -2940 -2468
rect -2906 -2502 -2873 -2468
rect -2974 -2702 -2873 -2502
rect -2974 -2736 -2940 -2702
rect -2906 -2736 -2873 -2702
rect -2974 -2770 -2873 -2736
rect -2974 -2804 -2940 -2770
rect -2906 -2804 -2873 -2770
rect -2974 -2838 -2873 -2804
rect -2811 -2417 -2393 -2393
rect -2811 -2451 -2787 -2417
rect -2753 -2451 -2719 -2417
rect -2685 -2451 -2519 -2417
rect -2485 -2451 -2451 -2417
rect -2417 -2451 -2393 -2417
rect -2811 -2465 -2393 -2451
rect -2811 -2485 -2739 -2465
rect -2811 -2519 -2787 -2485
rect -2753 -2519 -2739 -2485
rect -2811 -2685 -2739 -2519
rect -2465 -2485 -2393 -2465
rect -2465 -2519 -2451 -2485
rect -2417 -2519 -2393 -2485
rect -2681 -2537 -2523 -2523
rect -2681 -2571 -2667 -2537
rect -2633 -2551 -2571 -2537
rect -2537 -2571 -2523 -2537
rect -2681 -2633 -2653 -2571
rect -2551 -2633 -2523 -2571
rect -2681 -2667 -2667 -2633
rect -2633 -2667 -2571 -2653
rect -2537 -2667 -2523 -2633
rect -2681 -2681 -2523 -2667
rect -2811 -2719 -2787 -2685
rect -2753 -2719 -2739 -2685
rect -2811 -2739 -2739 -2719
rect -2465 -2685 -2393 -2519
rect -2465 -2719 -2451 -2685
rect -2417 -2719 -2393 -2685
rect -2465 -2739 -2393 -2719
rect -2811 -2753 -2393 -2739
rect -2811 -2787 -2787 -2753
rect -2753 -2787 -2719 -2753
rect -2685 -2787 -2519 -2753
rect -2485 -2787 -2451 -2753
rect -2417 -2787 -2393 -2753
rect -2811 -2811 -2393 -2787
rect -2331 -2400 -2230 -2366
rect -2331 -2434 -2298 -2400
rect -2264 -2434 -2230 -2400
rect -2331 -2468 -2230 -2434
rect -2331 -2502 -2298 -2468
rect -2264 -2502 -2230 -2468
rect -2331 -2702 -2230 -2502
rect -2331 -2736 -2298 -2702
rect -2264 -2736 -2230 -2702
rect -2331 -2770 -2230 -2736
rect -2331 -2804 -2298 -2770
rect -2264 -2804 -2230 -2770
rect -2974 -2872 -2940 -2838
rect -2906 -2872 -2873 -2838
rect -2974 -2873 -2873 -2872
rect -2331 -2838 -2230 -2804
rect -2331 -2872 -2298 -2838
rect -2264 -2872 -2230 -2838
rect -2331 -2873 -2230 -2872
rect -2974 -2906 -2230 -2873
rect -2974 -2940 -2940 -2906
rect -2906 -2940 -2872 -2906
rect -2838 -2940 -2804 -2906
rect -2770 -2940 -2736 -2906
rect -2702 -2940 -2502 -2906
rect -2468 -2940 -2434 -2906
rect -2400 -2940 -2366 -2906
rect -2332 -2940 -2298 -2906
rect -2264 -2940 -2230 -2906
rect -2974 -2974 -2230 -2940
rect -1974 -2264 -1230 -2230
rect -1974 -2298 -1940 -2264
rect -1906 -2298 -1872 -2264
rect -1838 -2298 -1804 -2264
rect -1770 -2298 -1736 -2264
rect -1702 -2298 -1502 -2264
rect -1468 -2298 -1434 -2264
rect -1400 -2298 -1366 -2264
rect -1332 -2298 -1298 -2264
rect -1264 -2298 -1230 -2264
rect -1974 -2331 -1230 -2298
rect -1974 -2332 -1873 -2331
rect -1974 -2366 -1940 -2332
rect -1906 -2366 -1873 -2332
rect -1974 -2400 -1873 -2366
rect -1331 -2332 -1230 -2331
rect -1331 -2366 -1298 -2332
rect -1264 -2366 -1230 -2332
rect -1974 -2434 -1940 -2400
rect -1906 -2434 -1873 -2400
rect -1974 -2468 -1873 -2434
rect -1974 -2502 -1940 -2468
rect -1906 -2502 -1873 -2468
rect -1974 -2702 -1873 -2502
rect -1974 -2736 -1940 -2702
rect -1906 -2736 -1873 -2702
rect -1974 -2770 -1873 -2736
rect -1974 -2804 -1940 -2770
rect -1906 -2804 -1873 -2770
rect -1974 -2838 -1873 -2804
rect -1811 -2417 -1393 -2393
rect -1811 -2451 -1787 -2417
rect -1753 -2451 -1719 -2417
rect -1685 -2451 -1519 -2417
rect -1485 -2451 -1451 -2417
rect -1417 -2451 -1393 -2417
rect -1811 -2465 -1393 -2451
rect -1811 -2485 -1739 -2465
rect -1811 -2519 -1787 -2485
rect -1753 -2519 -1739 -2485
rect -1811 -2685 -1739 -2519
rect -1465 -2485 -1393 -2465
rect -1465 -2519 -1451 -2485
rect -1417 -2519 -1393 -2485
rect -1681 -2537 -1523 -2523
rect -1681 -2571 -1667 -2537
rect -1633 -2551 -1571 -2537
rect -1537 -2571 -1523 -2537
rect -1681 -2633 -1653 -2571
rect -1551 -2633 -1523 -2571
rect -1681 -2667 -1667 -2633
rect -1633 -2667 -1571 -2653
rect -1537 -2667 -1523 -2633
rect -1681 -2681 -1523 -2667
rect -1811 -2719 -1787 -2685
rect -1753 -2719 -1739 -2685
rect -1811 -2739 -1739 -2719
rect -1465 -2685 -1393 -2519
rect -1465 -2719 -1451 -2685
rect -1417 -2719 -1393 -2685
rect -1465 -2739 -1393 -2719
rect -1811 -2753 -1393 -2739
rect -1811 -2787 -1787 -2753
rect -1753 -2787 -1719 -2753
rect -1685 -2787 -1519 -2753
rect -1485 -2787 -1451 -2753
rect -1417 -2787 -1393 -2753
rect -1811 -2811 -1393 -2787
rect -1331 -2400 -1230 -2366
rect -1331 -2434 -1298 -2400
rect -1264 -2434 -1230 -2400
rect -1331 -2468 -1230 -2434
rect -1331 -2502 -1298 -2468
rect -1264 -2502 -1230 -2468
rect -1331 -2702 -1230 -2502
rect -1331 -2736 -1298 -2702
rect -1264 -2736 -1230 -2702
rect -1331 -2770 -1230 -2736
rect -1331 -2804 -1298 -2770
rect -1264 -2804 -1230 -2770
rect -1974 -2872 -1940 -2838
rect -1906 -2872 -1873 -2838
rect -1974 -2873 -1873 -2872
rect -1331 -2838 -1230 -2804
rect -1331 -2872 -1298 -2838
rect -1264 -2872 -1230 -2838
rect -1331 -2873 -1230 -2872
rect -1974 -2906 -1230 -2873
rect -1974 -2940 -1940 -2906
rect -1906 -2940 -1872 -2906
rect -1838 -2940 -1804 -2906
rect -1770 -2940 -1736 -2906
rect -1702 -2940 -1502 -2906
rect -1468 -2940 -1434 -2906
rect -1400 -2940 -1366 -2906
rect -1332 -2940 -1298 -2906
rect -1264 -2940 -1230 -2906
rect -1974 -2974 -1230 -2940
rect -974 -2264 -230 -2230
rect -974 -2298 -940 -2264
rect -906 -2298 -872 -2264
rect -838 -2298 -804 -2264
rect -770 -2298 -736 -2264
rect -702 -2298 -502 -2264
rect -468 -2298 -434 -2264
rect -400 -2298 -366 -2264
rect -332 -2298 -298 -2264
rect -264 -2298 -230 -2264
rect -974 -2331 -230 -2298
rect -974 -2332 -873 -2331
rect -974 -2366 -940 -2332
rect -906 -2366 -873 -2332
rect -974 -2400 -873 -2366
rect -331 -2332 -230 -2331
rect -331 -2366 -298 -2332
rect -264 -2366 -230 -2332
rect -974 -2434 -940 -2400
rect -906 -2434 -873 -2400
rect -974 -2468 -873 -2434
rect -974 -2502 -940 -2468
rect -906 -2502 -873 -2468
rect -974 -2702 -873 -2502
rect -974 -2736 -940 -2702
rect -906 -2736 -873 -2702
rect -974 -2770 -873 -2736
rect -974 -2804 -940 -2770
rect -906 -2804 -873 -2770
rect -974 -2838 -873 -2804
rect -811 -2417 -393 -2393
rect -811 -2451 -787 -2417
rect -753 -2451 -719 -2417
rect -685 -2451 -519 -2417
rect -485 -2451 -451 -2417
rect -417 -2451 -393 -2417
rect -811 -2465 -393 -2451
rect -811 -2485 -739 -2465
rect -811 -2519 -787 -2485
rect -753 -2519 -739 -2485
rect -811 -2685 -739 -2519
rect -465 -2485 -393 -2465
rect -465 -2519 -451 -2485
rect -417 -2519 -393 -2485
rect -681 -2537 -523 -2523
rect -681 -2571 -667 -2537
rect -633 -2551 -571 -2537
rect -537 -2571 -523 -2537
rect -681 -2633 -653 -2571
rect -551 -2633 -523 -2571
rect -681 -2667 -667 -2633
rect -633 -2667 -571 -2653
rect -537 -2667 -523 -2633
rect -681 -2681 -523 -2667
rect -811 -2719 -787 -2685
rect -753 -2719 -739 -2685
rect -811 -2739 -739 -2719
rect -465 -2685 -393 -2519
rect -465 -2719 -451 -2685
rect -417 -2719 -393 -2685
rect -465 -2739 -393 -2719
rect -811 -2753 -393 -2739
rect -811 -2787 -787 -2753
rect -753 -2787 -719 -2753
rect -685 -2787 -519 -2753
rect -485 -2787 -451 -2753
rect -417 -2787 -393 -2753
rect -811 -2811 -393 -2787
rect -331 -2400 -230 -2366
rect -331 -2434 -298 -2400
rect -264 -2434 -230 -2400
rect -331 -2468 -230 -2434
rect -331 -2502 -298 -2468
rect -264 -2502 -230 -2468
rect -331 -2702 -230 -2502
rect -331 -2736 -298 -2702
rect -264 -2736 -230 -2702
rect -331 -2770 -230 -2736
rect -331 -2804 -298 -2770
rect -264 -2804 -230 -2770
rect -974 -2872 -940 -2838
rect -906 -2872 -873 -2838
rect -974 -2873 -873 -2872
rect -331 -2838 -230 -2804
rect -331 -2872 -298 -2838
rect -264 -2872 -230 -2838
rect -331 -2873 -230 -2872
rect -974 -2906 -230 -2873
rect -974 -2940 -940 -2906
rect -906 -2940 -872 -2906
rect -838 -2940 -804 -2906
rect -770 -2940 -736 -2906
rect -702 -2940 -502 -2906
rect -468 -2940 -434 -2906
rect -400 -2940 -366 -2906
rect -332 -2940 -298 -2906
rect -264 -2940 -230 -2906
rect -974 -2974 -230 -2940
rect 26 -2264 770 -2230
rect 26 -2298 60 -2264
rect 94 -2298 128 -2264
rect 162 -2298 196 -2264
rect 230 -2298 264 -2264
rect 298 -2298 498 -2264
rect 532 -2298 566 -2264
rect 600 -2298 634 -2264
rect 668 -2298 702 -2264
rect 736 -2298 770 -2264
rect 26 -2331 770 -2298
rect 26 -2332 127 -2331
rect 26 -2366 60 -2332
rect 94 -2366 127 -2332
rect 26 -2400 127 -2366
rect 669 -2332 770 -2331
rect 669 -2366 702 -2332
rect 736 -2366 770 -2332
rect 26 -2434 60 -2400
rect 94 -2434 127 -2400
rect 26 -2468 127 -2434
rect 26 -2502 60 -2468
rect 94 -2502 127 -2468
rect 26 -2702 127 -2502
rect 26 -2736 60 -2702
rect 94 -2736 127 -2702
rect 26 -2770 127 -2736
rect 26 -2804 60 -2770
rect 94 -2804 127 -2770
rect 26 -2838 127 -2804
rect 189 -2417 607 -2393
rect 189 -2451 213 -2417
rect 247 -2451 281 -2417
rect 315 -2451 481 -2417
rect 515 -2451 549 -2417
rect 583 -2451 607 -2417
rect 189 -2465 607 -2451
rect 189 -2485 261 -2465
rect 189 -2519 213 -2485
rect 247 -2519 261 -2485
rect 189 -2685 261 -2519
rect 535 -2485 607 -2465
rect 535 -2519 549 -2485
rect 583 -2519 607 -2485
rect 319 -2537 477 -2523
rect 319 -2571 333 -2537
rect 367 -2551 429 -2537
rect 463 -2571 477 -2537
rect 319 -2633 347 -2571
rect 449 -2633 477 -2571
rect 319 -2667 333 -2633
rect 367 -2667 429 -2653
rect 463 -2667 477 -2633
rect 319 -2681 477 -2667
rect 189 -2719 213 -2685
rect 247 -2719 261 -2685
rect 189 -2739 261 -2719
rect 535 -2685 607 -2519
rect 535 -2719 549 -2685
rect 583 -2719 607 -2685
rect 535 -2739 607 -2719
rect 189 -2753 607 -2739
rect 189 -2787 213 -2753
rect 247 -2787 281 -2753
rect 315 -2787 481 -2753
rect 515 -2787 549 -2753
rect 583 -2787 607 -2753
rect 189 -2811 607 -2787
rect 669 -2400 770 -2366
rect 669 -2434 702 -2400
rect 736 -2434 770 -2400
rect 669 -2468 770 -2434
rect 669 -2502 702 -2468
rect 736 -2502 770 -2468
rect 669 -2702 770 -2502
rect 669 -2736 702 -2702
rect 736 -2736 770 -2702
rect 669 -2770 770 -2736
rect 669 -2804 702 -2770
rect 736 -2804 770 -2770
rect 26 -2872 60 -2838
rect 94 -2872 127 -2838
rect 26 -2873 127 -2872
rect 669 -2838 770 -2804
rect 669 -2872 702 -2838
rect 736 -2872 770 -2838
rect 669 -2873 770 -2872
rect 26 -2906 770 -2873
rect 26 -2940 60 -2906
rect 94 -2940 128 -2906
rect 162 -2940 196 -2906
rect 230 -2940 264 -2906
rect 298 -2940 498 -2906
rect 532 -2940 566 -2906
rect 600 -2940 634 -2906
rect 668 -2940 702 -2906
rect 736 -2940 770 -2906
rect 26 -2974 770 -2940
rect 1026 -2264 1770 -2230
rect 1026 -2298 1060 -2264
rect 1094 -2298 1128 -2264
rect 1162 -2298 1196 -2264
rect 1230 -2298 1264 -2264
rect 1298 -2298 1498 -2264
rect 1532 -2298 1566 -2264
rect 1600 -2298 1634 -2264
rect 1668 -2298 1702 -2264
rect 1736 -2298 1770 -2264
rect 1026 -2331 1770 -2298
rect 1026 -2332 1127 -2331
rect 1026 -2366 1060 -2332
rect 1094 -2366 1127 -2332
rect 1026 -2400 1127 -2366
rect 1669 -2332 1770 -2331
rect 1669 -2366 1702 -2332
rect 1736 -2366 1770 -2332
rect 1026 -2434 1060 -2400
rect 1094 -2434 1127 -2400
rect 1026 -2468 1127 -2434
rect 1026 -2502 1060 -2468
rect 1094 -2502 1127 -2468
rect 1026 -2702 1127 -2502
rect 1026 -2736 1060 -2702
rect 1094 -2736 1127 -2702
rect 1026 -2770 1127 -2736
rect 1026 -2804 1060 -2770
rect 1094 -2804 1127 -2770
rect 1026 -2838 1127 -2804
rect 1189 -2417 1607 -2393
rect 1189 -2451 1213 -2417
rect 1247 -2451 1281 -2417
rect 1315 -2451 1481 -2417
rect 1515 -2451 1549 -2417
rect 1583 -2451 1607 -2417
rect 1189 -2465 1607 -2451
rect 1189 -2485 1261 -2465
rect 1189 -2519 1213 -2485
rect 1247 -2519 1261 -2485
rect 1189 -2685 1261 -2519
rect 1535 -2485 1607 -2465
rect 1535 -2519 1549 -2485
rect 1583 -2519 1607 -2485
rect 1319 -2537 1477 -2523
rect 1319 -2571 1333 -2537
rect 1367 -2551 1429 -2537
rect 1463 -2571 1477 -2537
rect 1319 -2633 1347 -2571
rect 1449 -2633 1477 -2571
rect 1319 -2667 1333 -2633
rect 1367 -2667 1429 -2653
rect 1463 -2667 1477 -2633
rect 1319 -2681 1477 -2667
rect 1189 -2719 1213 -2685
rect 1247 -2719 1261 -2685
rect 1189 -2739 1261 -2719
rect 1535 -2685 1607 -2519
rect 1535 -2719 1549 -2685
rect 1583 -2719 1607 -2685
rect 1535 -2739 1607 -2719
rect 1189 -2753 1607 -2739
rect 1189 -2787 1213 -2753
rect 1247 -2787 1281 -2753
rect 1315 -2787 1481 -2753
rect 1515 -2787 1549 -2753
rect 1583 -2787 1607 -2753
rect 1189 -2811 1607 -2787
rect 1669 -2400 1770 -2366
rect 1669 -2434 1702 -2400
rect 1736 -2434 1770 -2400
rect 1669 -2468 1770 -2434
rect 1669 -2502 1702 -2468
rect 1736 -2502 1770 -2468
rect 1669 -2702 1770 -2502
rect 1669 -2736 1702 -2702
rect 1736 -2736 1770 -2702
rect 1669 -2770 1770 -2736
rect 1669 -2804 1702 -2770
rect 1736 -2804 1770 -2770
rect 1026 -2872 1060 -2838
rect 1094 -2872 1127 -2838
rect 1026 -2873 1127 -2872
rect 1669 -2838 1770 -2804
rect 1669 -2872 1702 -2838
rect 1736 -2872 1770 -2838
rect 1669 -2873 1770 -2872
rect 1026 -2906 1770 -2873
rect 1026 -2940 1060 -2906
rect 1094 -2940 1128 -2906
rect 1162 -2940 1196 -2906
rect 1230 -2940 1264 -2906
rect 1298 -2940 1498 -2906
rect 1532 -2940 1566 -2906
rect 1600 -2940 1634 -2906
rect 1668 -2940 1702 -2906
rect 1736 -2940 1770 -2906
rect 1026 -2974 1770 -2940
<< viali >>
rect -3667 1449 -3633 1463
rect -3571 1449 -3537 1463
rect -3667 1429 -3653 1449
rect -3653 1429 -3633 1449
rect -3571 1429 -3551 1449
rect -3551 1429 -3537 1449
rect -3667 1347 -3653 1367
rect -3653 1347 -3633 1367
rect -3571 1347 -3551 1367
rect -3551 1347 -3537 1367
rect -3667 1333 -3633 1347
rect -3571 1333 -3537 1347
rect -2667 1449 -2633 1463
rect -2571 1449 -2537 1463
rect -2667 1429 -2653 1449
rect -2653 1429 -2633 1449
rect -2571 1429 -2551 1449
rect -2551 1429 -2537 1449
rect -2667 1347 -2653 1367
rect -2653 1347 -2633 1367
rect -2571 1347 -2551 1367
rect -2551 1347 -2537 1367
rect -2667 1333 -2633 1347
rect -2571 1333 -2537 1347
rect -1667 1449 -1633 1463
rect -1571 1449 -1537 1463
rect -1667 1429 -1653 1449
rect -1653 1429 -1633 1449
rect -1571 1429 -1551 1449
rect -1551 1429 -1537 1449
rect -1667 1347 -1653 1367
rect -1653 1347 -1633 1367
rect -1571 1347 -1551 1367
rect -1551 1347 -1537 1367
rect -1667 1333 -1633 1347
rect -1571 1333 -1537 1347
rect -667 1449 -633 1463
rect -571 1449 -537 1463
rect -667 1429 -653 1449
rect -653 1429 -633 1449
rect -571 1429 -551 1449
rect -551 1429 -537 1449
rect -667 1347 -653 1367
rect -653 1347 -633 1367
rect -571 1347 -551 1367
rect -551 1347 -537 1367
rect -667 1333 -633 1347
rect -571 1333 -537 1347
rect 333 1449 367 1463
rect 429 1449 463 1463
rect 333 1429 347 1449
rect 347 1429 367 1449
rect 429 1429 449 1449
rect 449 1429 463 1449
rect 333 1347 347 1367
rect 347 1347 367 1367
rect 429 1347 449 1367
rect 449 1347 463 1367
rect 333 1333 367 1347
rect 429 1333 463 1347
rect 1333 1449 1367 1463
rect 1429 1449 1463 1463
rect 1333 1429 1347 1449
rect 1347 1429 1367 1449
rect 1429 1429 1449 1449
rect 1449 1429 1463 1449
rect 1333 1347 1347 1367
rect 1347 1347 1367 1367
rect 1429 1347 1449 1367
rect 1449 1347 1463 1367
rect 1333 1333 1367 1347
rect 1429 1333 1463 1347
rect -3667 449 -3633 463
rect -3571 449 -3537 463
rect -3667 429 -3653 449
rect -3653 429 -3633 449
rect -3571 429 -3551 449
rect -3551 429 -3537 449
rect -3667 347 -3653 367
rect -3653 347 -3633 367
rect -3571 347 -3551 367
rect -3551 347 -3537 367
rect -3667 333 -3633 347
rect -3571 333 -3537 347
rect -2667 449 -2633 463
rect -2571 449 -2537 463
rect -2667 429 -2653 449
rect -2653 429 -2633 449
rect -2571 429 -2551 449
rect -2551 429 -2537 449
rect -2667 347 -2653 367
rect -2653 347 -2633 367
rect -2571 347 -2551 367
rect -2551 347 -2537 367
rect -2667 333 -2633 347
rect -2571 333 -2537 347
rect -1667 449 -1633 463
rect -1571 449 -1537 463
rect -1667 429 -1653 449
rect -1653 429 -1633 449
rect -1571 429 -1551 449
rect -1551 429 -1537 449
rect -1667 347 -1653 367
rect -1653 347 -1633 367
rect -1571 347 -1551 367
rect -1551 347 -1537 367
rect -1667 333 -1633 347
rect -1571 333 -1537 347
rect -667 449 -633 463
rect -571 449 -537 463
rect -667 429 -653 449
rect -653 429 -633 449
rect -571 429 -551 449
rect -551 429 -537 449
rect -667 347 -653 367
rect -653 347 -633 367
rect -571 347 -551 367
rect -551 347 -537 367
rect -667 333 -633 347
rect -571 333 -537 347
rect 333 449 367 463
rect 429 449 463 463
rect 333 429 347 449
rect 347 429 367 449
rect 429 429 449 449
rect 449 429 463 449
rect 333 347 347 367
rect 347 347 367 367
rect 429 347 449 367
rect 449 347 463 367
rect 333 333 367 347
rect 429 333 463 347
rect 1333 449 1367 463
rect 1429 449 1463 463
rect 1333 429 1347 449
rect 1347 429 1367 449
rect 1429 429 1449 449
rect 1449 429 1463 449
rect 1333 347 1347 367
rect 1347 347 1367 367
rect 1429 347 1449 367
rect 1449 347 1463 367
rect 1333 333 1367 347
rect 1429 333 1463 347
rect -3667 -551 -3633 -537
rect -3571 -551 -3537 -537
rect -3667 -571 -3653 -551
rect -3653 -571 -3633 -551
rect -3571 -571 -3551 -551
rect -3551 -571 -3537 -551
rect -3667 -653 -3653 -633
rect -3653 -653 -3633 -633
rect -3571 -653 -3551 -633
rect -3551 -653 -3537 -633
rect -3667 -667 -3633 -653
rect -3571 -667 -3537 -653
rect -2667 -551 -2633 -537
rect -2571 -551 -2537 -537
rect -2667 -571 -2653 -551
rect -2653 -571 -2633 -551
rect -2571 -571 -2551 -551
rect -2551 -571 -2537 -551
rect -2667 -653 -2653 -633
rect -2653 -653 -2633 -633
rect -2571 -653 -2551 -633
rect -2551 -653 -2537 -633
rect -2667 -667 -2633 -653
rect -2571 -667 -2537 -653
rect -1667 -551 -1633 -537
rect -1571 -551 -1537 -537
rect -1667 -571 -1653 -551
rect -1653 -571 -1633 -551
rect -1571 -571 -1551 -551
rect -1551 -571 -1537 -551
rect -1667 -653 -1653 -633
rect -1653 -653 -1633 -633
rect -1571 -653 -1551 -633
rect -1551 -653 -1537 -633
rect -1667 -667 -1633 -653
rect -1571 -667 -1537 -653
rect -667 -551 -633 -537
rect -571 -551 -537 -537
rect -667 -571 -653 -551
rect -653 -571 -633 -551
rect -571 -571 -551 -551
rect -551 -571 -537 -551
rect -667 -653 -653 -633
rect -653 -653 -633 -633
rect -571 -653 -551 -633
rect -551 -653 -537 -633
rect -667 -667 -633 -653
rect -571 -667 -537 -653
rect 333 -551 367 -537
rect 429 -551 463 -537
rect 333 -571 347 -551
rect 347 -571 367 -551
rect 429 -571 449 -551
rect 449 -571 463 -551
rect 333 -653 347 -633
rect 347 -653 367 -633
rect 429 -653 449 -633
rect 449 -653 463 -633
rect 333 -667 367 -653
rect 429 -667 463 -653
rect 1333 -551 1367 -537
rect 1429 -551 1463 -537
rect 1333 -571 1347 -551
rect 1347 -571 1367 -551
rect 1429 -571 1449 -551
rect 1449 -571 1463 -551
rect 1333 -653 1347 -633
rect 1347 -653 1367 -633
rect 1429 -653 1449 -633
rect 1449 -653 1463 -633
rect 1333 -667 1367 -653
rect 1429 -667 1463 -653
rect -3667 -1551 -3633 -1537
rect -3571 -1551 -3537 -1537
rect -3667 -1571 -3653 -1551
rect -3653 -1571 -3633 -1551
rect -3571 -1571 -3551 -1551
rect -3551 -1571 -3537 -1551
rect -3667 -1653 -3653 -1633
rect -3653 -1653 -3633 -1633
rect -3571 -1653 -3551 -1633
rect -3551 -1653 -3537 -1633
rect -3667 -1667 -3633 -1653
rect -3571 -1667 -3537 -1653
rect -2667 -1551 -2633 -1537
rect -2571 -1551 -2537 -1537
rect -2667 -1571 -2653 -1551
rect -2653 -1571 -2633 -1551
rect -2571 -1571 -2551 -1551
rect -2551 -1571 -2537 -1551
rect -2667 -1653 -2653 -1633
rect -2653 -1653 -2633 -1633
rect -2571 -1653 -2551 -1633
rect -2551 -1653 -2537 -1633
rect -2667 -1667 -2633 -1653
rect -2571 -1667 -2537 -1653
rect -1667 -1551 -1633 -1537
rect -1571 -1551 -1537 -1537
rect -1667 -1571 -1653 -1551
rect -1653 -1571 -1633 -1551
rect -1571 -1571 -1551 -1551
rect -1551 -1571 -1537 -1551
rect -1667 -1653 -1653 -1633
rect -1653 -1653 -1633 -1633
rect -1571 -1653 -1551 -1633
rect -1551 -1653 -1537 -1633
rect -1667 -1667 -1633 -1653
rect -1571 -1667 -1537 -1653
rect -667 -1551 -633 -1537
rect -571 -1551 -537 -1537
rect -667 -1571 -653 -1551
rect -653 -1571 -633 -1551
rect -571 -1571 -551 -1551
rect -551 -1571 -537 -1551
rect -667 -1653 -653 -1633
rect -653 -1653 -633 -1633
rect -571 -1653 -551 -1633
rect -551 -1653 -537 -1633
rect -667 -1667 -633 -1653
rect -571 -1667 -537 -1653
rect 550 -1417 590 -1410
rect 550 -1450 583 -1417
rect 583 -1450 590 -1417
rect 333 -1551 367 -1537
rect 429 -1551 463 -1537
rect 333 -1571 347 -1551
rect 347 -1571 367 -1551
rect 429 -1571 449 -1551
rect 449 -1571 463 -1551
rect 333 -1653 347 -1633
rect 347 -1653 367 -1633
rect 429 -1653 449 -1633
rect 449 -1653 463 -1633
rect 333 -1667 367 -1653
rect 429 -1667 463 -1653
rect 700 -1906 740 -1900
rect 700 -1940 702 -1906
rect 702 -1940 736 -1906
rect 736 -1940 740 -1906
rect 2250 -1320 2300 -920
rect 1333 -1551 1367 -1537
rect 1429 -1551 1463 -1537
rect 1333 -1571 1347 -1551
rect 1347 -1571 1367 -1551
rect 1429 -1571 1449 -1551
rect 1449 -1571 1463 -1551
rect 1333 -1653 1347 -1633
rect 1347 -1653 1367 -1633
rect 1429 -1653 1449 -1633
rect 1449 -1653 1463 -1633
rect 1333 -1667 1367 -1653
rect 1429 -1667 1463 -1653
rect -3667 -2551 -3633 -2537
rect -3571 -2551 -3537 -2537
rect -3667 -2571 -3653 -2551
rect -3653 -2571 -3633 -2551
rect -3571 -2571 -3551 -2551
rect -3551 -2571 -3537 -2551
rect -3667 -2653 -3653 -2633
rect -3653 -2653 -3633 -2633
rect -3571 -2653 -3551 -2633
rect -3551 -2653 -3537 -2633
rect -3667 -2667 -3633 -2653
rect -3571 -2667 -3537 -2653
rect -2667 -2551 -2633 -2537
rect -2571 -2551 -2537 -2537
rect -2667 -2571 -2653 -2551
rect -2653 -2571 -2633 -2551
rect -2571 -2571 -2551 -2551
rect -2551 -2571 -2537 -2551
rect -2667 -2653 -2653 -2633
rect -2653 -2653 -2633 -2633
rect -2571 -2653 -2551 -2633
rect -2551 -2653 -2537 -2633
rect -2667 -2667 -2633 -2653
rect -2571 -2667 -2537 -2653
rect -1667 -2551 -1633 -2537
rect -1571 -2551 -1537 -2537
rect -1667 -2571 -1653 -2551
rect -1653 -2571 -1633 -2551
rect -1571 -2571 -1551 -2551
rect -1551 -2571 -1537 -2551
rect -1667 -2653 -1653 -2633
rect -1653 -2653 -1633 -2633
rect -1571 -2653 -1551 -2633
rect -1551 -2653 -1537 -2633
rect -1667 -2667 -1633 -2653
rect -1571 -2667 -1537 -2653
rect -667 -2551 -633 -2537
rect -571 -2551 -537 -2537
rect -667 -2571 -653 -2551
rect -653 -2571 -633 -2551
rect -571 -2571 -551 -2551
rect -551 -2571 -537 -2551
rect -667 -2653 -653 -2633
rect -653 -2653 -633 -2633
rect -571 -2653 -551 -2633
rect -551 -2653 -537 -2633
rect -667 -2667 -633 -2653
rect -571 -2667 -537 -2653
rect 333 -2551 367 -2537
rect 429 -2551 463 -2537
rect 333 -2571 347 -2551
rect 347 -2571 367 -2551
rect 429 -2571 449 -2551
rect 449 -2571 463 -2551
rect 333 -2653 347 -2633
rect 347 -2653 367 -2633
rect 429 -2653 449 -2633
rect 449 -2653 463 -2633
rect 333 -2667 367 -2653
rect 429 -2667 463 -2653
rect 1333 -2551 1367 -2537
rect 1429 -2551 1463 -2537
rect 1333 -2571 1347 -2551
rect 1347 -2571 1367 -2551
rect 1429 -2571 1449 -2551
rect 1449 -2571 1463 -2551
rect 1333 -2653 1347 -2633
rect 1347 -2653 1367 -2633
rect 1429 -2653 1449 -2633
rect 1449 -2653 1463 -2633
rect 1333 -2667 1367 -2653
rect 1429 -2667 1463 -2653
rect 2250 -2460 2300 -2060
rect -810 -3360 -410 -3310
rect -110 -3360 290 -3310
<< metal1 >>
rect -3685 1463 -3519 1481
rect -3685 1429 -3667 1463
rect -3633 1429 -3571 1463
rect -3537 1429 -3519 1463
rect -3685 1367 -3519 1429
rect -3685 1333 -3667 1367
rect -3633 1333 -3571 1367
rect -3537 1333 -3519 1367
rect -3685 1315 -3519 1333
rect -2685 1463 -2519 1481
rect -2685 1429 -2667 1463
rect -2633 1429 -2571 1463
rect -2537 1429 -2519 1463
rect -2685 1367 -2519 1429
rect -2685 1333 -2667 1367
rect -2633 1333 -2571 1367
rect -2537 1333 -2519 1367
rect -2685 1315 -2519 1333
rect -1685 1463 -1519 1481
rect -1685 1429 -1667 1463
rect -1633 1429 -1571 1463
rect -1537 1429 -1519 1463
rect -1685 1367 -1519 1429
rect -1685 1333 -1667 1367
rect -1633 1333 -1571 1367
rect -1537 1333 -1519 1367
rect -1685 1315 -1519 1333
rect -685 1463 -519 1481
rect -685 1429 -667 1463
rect -633 1429 -571 1463
rect -537 1429 -519 1463
rect -685 1367 -519 1429
rect -685 1333 -667 1367
rect -633 1333 -571 1367
rect -537 1333 -519 1367
rect -685 1315 -519 1333
rect 315 1463 481 1481
rect 315 1429 333 1463
rect 367 1429 429 1463
rect 463 1429 481 1463
rect 315 1367 481 1429
rect 315 1333 333 1367
rect 367 1333 429 1367
rect 463 1333 481 1367
rect 315 1315 481 1333
rect 1315 1463 1481 1481
rect 1315 1429 1333 1463
rect 1367 1429 1429 1463
rect 1463 1429 1481 1463
rect 1315 1367 1481 1429
rect 1315 1333 1333 1367
rect 1367 1333 1429 1367
rect 1463 1333 1481 1367
rect 1315 1315 1481 1333
rect -3685 463 -3519 481
rect -3685 429 -3667 463
rect -3633 429 -3571 463
rect -3537 429 -3519 463
rect -3685 367 -3519 429
rect -3685 333 -3667 367
rect -3633 333 -3571 367
rect -3537 333 -3519 367
rect -3685 315 -3519 333
rect -2685 480 -2519 481
rect -1685 480 -1519 481
rect -685 480 -519 481
rect -2685 463 -519 480
rect -2685 429 -2667 463
rect -2633 429 -2571 463
rect -2537 429 -1667 463
rect -1633 429 -1571 463
rect -1537 429 -667 463
rect -633 429 -571 463
rect -537 429 -519 463
rect -2685 367 -519 429
rect -2685 333 -2667 367
rect -2633 333 -2571 367
rect -2537 333 -1667 367
rect -1633 333 -1571 367
rect -1537 333 -667 367
rect -633 333 -571 367
rect -537 333 -519 367
rect -2685 320 -519 333
rect -2685 315 -2519 320
rect -1685 315 -1519 320
rect -685 315 -519 320
rect 315 463 481 481
rect 315 429 333 463
rect 367 429 429 463
rect 463 429 481 463
rect 315 367 481 429
rect 315 333 333 367
rect 367 333 429 367
rect 463 333 481 367
rect 315 315 481 333
rect 1315 463 1481 481
rect 1315 429 1333 463
rect 1367 429 1429 463
rect 1463 429 1481 463
rect 1315 367 1481 429
rect 1315 333 1333 367
rect 1367 333 1429 367
rect 1463 333 1481 367
rect 1315 315 1481 333
rect -2680 -519 -2530 315
rect -1680 -519 -1530 315
rect -680 -519 -520 315
rect -3685 -537 -3519 -519
rect -3685 -571 -3667 -537
rect -3633 -571 -3571 -537
rect -3537 -571 -3519 -537
rect -3685 -633 -3519 -571
rect -3685 -667 -3667 -633
rect -3633 -667 -3571 -633
rect -3537 -667 -3519 -633
rect -3685 -685 -3519 -667
rect -2685 -520 -2519 -519
rect -1685 -520 -1519 -519
rect -685 -520 -519 -519
rect -2685 -537 -519 -520
rect -2685 -571 -2667 -537
rect -2633 -571 -2571 -537
rect -2537 -571 -1667 -537
rect -1633 -571 -1571 -537
rect -1537 -571 -667 -537
rect -633 -571 -571 -537
rect -537 -571 -519 -537
rect -2685 -633 -519 -571
rect -2685 -667 -2667 -633
rect -2633 -667 -2571 -633
rect -2537 -667 -1667 -633
rect -1633 -667 -1571 -633
rect -1537 -667 -667 -633
rect -633 -667 -571 -633
rect -537 -667 -519 -633
rect -2685 -680 -519 -667
rect -2685 -685 -2519 -680
rect -1685 -685 -1519 -680
rect -685 -685 -519 -680
rect 315 -537 481 -519
rect 315 -571 333 -537
rect 367 -571 429 -537
rect 463 -571 481 -537
rect 315 -633 481 -571
rect 315 -667 333 -633
rect 367 -667 429 -633
rect 463 -667 481 -633
rect 315 -685 481 -667
rect 1315 -537 1481 -519
rect 1315 -571 1333 -537
rect 1367 -571 1429 -537
rect 1463 -571 1481 -537
rect 1315 -633 1481 -571
rect 1315 -667 1333 -633
rect 1367 -667 1429 -633
rect 1463 -667 1481 -633
rect 1315 -685 1481 -667
rect -2680 -1510 -2530 -685
rect -1680 -1510 -1530 -685
rect 2240 -920 2310 -900
rect 2240 -1080 2250 -920
rect 870 -1120 2250 -1080
rect 870 -1400 910 -1120
rect 2240 -1320 2250 -1120
rect 2300 -1320 2310 -920
rect 2240 -1340 2310 -1320
rect 530 -1410 910 -1400
rect 530 -1450 550 -1410
rect 590 -1450 910 -1410
rect 530 -1470 910 -1450
rect -2680 -1519 -1520 -1510
rect -3685 -1537 -3519 -1519
rect -3685 -1571 -3667 -1537
rect -3633 -1571 -3571 -1537
rect -3537 -1571 -3519 -1537
rect -3685 -1633 -3519 -1571
rect -3685 -1667 -3667 -1633
rect -3633 -1667 -3571 -1633
rect -3537 -1667 -3519 -1633
rect -3685 -1685 -3519 -1667
rect -2685 -1537 -1519 -1519
rect -2685 -1571 -2667 -1537
rect -2633 -1571 -2571 -1537
rect -2537 -1571 -1667 -1537
rect -1633 -1571 -1571 -1537
rect -1537 -1571 -1519 -1537
rect -2685 -1633 -1519 -1571
rect -685 -1537 -519 -1519
rect -685 -1571 -667 -1537
rect -633 -1571 -571 -1537
rect -537 -1571 -519 -1537
rect -685 -1620 -519 -1571
rect -2685 -1667 -2667 -1633
rect -2633 -1667 -2571 -1633
rect -2537 -1667 -1667 -1633
rect -1633 -1667 -1571 -1633
rect -1537 -1667 -1519 -1633
rect -2685 -1680 -1519 -1667
rect -2685 -1685 -2519 -1680
rect -1685 -1685 -1519 -1680
rect -1130 -1633 -519 -1620
rect -1130 -1667 -667 -1633
rect -633 -1667 -571 -1633
rect -537 -1667 -519 -1633
rect -1130 -1680 -519 -1667
rect -3685 -2537 -3519 -2519
rect -3685 -2571 -3667 -2537
rect -3633 -2571 -3571 -2537
rect -3537 -2571 -3519 -2537
rect -3685 -2633 -3519 -2571
rect -3685 -2667 -3667 -2633
rect -3633 -2667 -3571 -2633
rect -3537 -2667 -3519 -2633
rect -3685 -2685 -3519 -2667
rect -2685 -2537 -2519 -2519
rect -2685 -2571 -2667 -2537
rect -2633 -2571 -2571 -2537
rect -2537 -2571 -2519 -2537
rect -2685 -2633 -2519 -2571
rect -2685 -2667 -2667 -2633
rect -2633 -2667 -2571 -2633
rect -2537 -2667 -2519 -2633
rect -2685 -2685 -2519 -2667
rect -1685 -2537 -1519 -2519
rect -1685 -2571 -1667 -2537
rect -1633 -2571 -1571 -2537
rect -1537 -2571 -1519 -2537
rect -1685 -2633 -1519 -2571
rect -1685 -2667 -1667 -2633
rect -1633 -2667 -1571 -2633
rect -1537 -2667 -1519 -2633
rect -1685 -2685 -1519 -2667
rect -1130 -3300 -1080 -1680
rect -685 -1685 -519 -1680
rect 315 -1537 481 -1519
rect 315 -1571 333 -1537
rect 367 -1571 429 -1537
rect 463 -1571 481 -1537
rect 315 -1633 481 -1571
rect 315 -1667 333 -1633
rect 367 -1667 429 -1633
rect 463 -1667 481 -1633
rect 315 -1685 481 -1667
rect 1315 -1537 1481 -1519
rect 1315 -1571 1333 -1537
rect 1367 -1571 1429 -1537
rect 1463 -1571 1481 -1537
rect 1315 -1633 1481 -1571
rect 1315 -1667 1333 -1633
rect 1367 -1667 1429 -1633
rect 1463 -1667 1481 -1633
rect 1315 -1685 1481 -1667
rect 670 -1900 910 -1870
rect 670 -1940 700 -1900
rect 740 -1940 910 -1900
rect 670 -1960 910 -1940
rect 870 -2100 910 -1960
rect 2240 -2060 2310 -2040
rect 2240 -2100 2250 -2060
rect 870 -2140 2250 -2100
rect 2240 -2460 2250 -2140
rect 2300 -2460 2310 -2060
rect 2240 -2480 2310 -2460
rect -685 -2537 -519 -2519
rect -685 -2571 -667 -2537
rect -633 -2571 -571 -2537
rect -537 -2571 -519 -2537
rect -685 -2633 -519 -2571
rect -685 -2667 -667 -2633
rect -633 -2667 -571 -2633
rect -537 -2667 -519 -2633
rect -685 -2685 -519 -2667
rect 315 -2537 481 -2519
rect 315 -2571 333 -2537
rect 367 -2571 429 -2537
rect 463 -2571 481 -2537
rect 315 -2633 481 -2571
rect 315 -2667 333 -2633
rect 367 -2667 429 -2633
rect 463 -2667 481 -2633
rect 315 -2685 481 -2667
rect 1315 -2537 1481 -2519
rect 1315 -2571 1333 -2537
rect 1367 -2571 1429 -2537
rect 1463 -2571 1481 -2537
rect 1315 -2633 1481 -2571
rect 1315 -2667 1333 -2633
rect 1367 -2667 1429 -2633
rect 1463 -2667 1481 -2633
rect 1315 -2685 1481 -2667
rect -1130 -3310 -390 -3300
rect -1130 -3360 -810 -3310
rect -410 -3360 -390 -3310
rect -1130 -3370 -390 -3360
rect -130 -3310 310 -3300
rect -130 -3360 -110 -3310
rect 290 -3360 310 -3310
rect -130 -3370 310 -3360
use p-res8x20k  p-res8x20k_0
timestamp 1620701388
transform 0 1 -140 -1 0 -3300
box 0 -1830 1180 1590
use p-res20k  p-res20k_0
timestamp 1620355008
transform 1 0 2240 0 1 -2040
box -200 -440 70 1140
<< end >>
