magic
tech sky130A
timestamp 1620435323
<< nwell >>
rect -120 370 85 610
<< nmos >>
rect 0 135 15 235
<< pmos >>
rect 0 390 15 590
<< ndiff >>
rect -50 220 0 235
rect -50 150 -35 220
rect -15 150 0 220
rect -50 135 0 150
rect 15 220 65 235
rect 15 150 30 220
rect 50 150 65 220
rect 15 135 65 150
<< pdiff >>
rect -50 575 0 590
rect -50 505 -35 575
rect -15 505 0 575
rect -50 475 0 505
rect -50 405 -35 475
rect -15 405 0 475
rect -50 390 0 405
rect 15 575 65 590
rect 15 505 30 575
rect 50 505 65 575
rect 15 475 65 505
rect 15 405 30 475
rect 50 405 65 475
rect 15 390 65 405
<< ndiffc >>
rect -35 150 -15 220
rect 30 150 50 220
<< pdiffc >>
rect -35 505 -15 575
rect -35 405 -15 475
rect 30 505 50 575
rect 30 405 50 475
<< psubdiff >>
rect -100 220 -50 235
rect -100 150 -85 220
rect -65 150 -50 220
rect -100 135 -50 150
<< nsubdiff >>
rect -100 575 -50 590
rect -100 505 -85 575
rect -65 505 -50 575
rect -100 475 -50 505
rect -100 405 -85 475
rect -65 405 -50 475
rect -100 390 -50 405
<< psubdiffcont >>
rect -85 150 -65 220
<< nsubdiffcont >>
rect -85 505 -65 575
rect -85 405 -65 475
<< poly >>
rect 0 590 15 605
rect 0 235 15 390
rect 0 120 15 135
rect -25 110 15 120
rect -25 90 -15 110
rect 5 90 15 110
rect -25 80 15 90
<< polycont >>
rect -15 90 5 110
<< locali >>
rect -95 575 -5 585
rect -95 505 -85 575
rect -65 505 -35 575
rect -15 505 -5 575
rect -95 475 -5 505
rect -95 405 -85 475
rect -65 405 -35 475
rect -15 405 -5 475
rect -95 395 -5 405
rect 20 575 60 585
rect 20 505 30 575
rect 50 505 60 575
rect 20 475 60 505
rect 20 405 30 475
rect 50 405 60 475
rect 20 395 60 405
rect 40 230 60 395
rect -95 220 -5 230
rect -95 150 -85 220
rect -65 150 -35 220
rect -15 150 -5 220
rect -95 140 -5 150
rect 20 220 60 230
rect 20 150 30 220
rect 50 150 60 220
rect 20 140 60 150
rect -25 110 15 120
rect -25 90 -15 110
rect 5 90 15 110
rect -25 80 15 90
rect 40 80 60 140
<< viali >>
rect -85 505 -65 575
rect -35 505 -15 575
rect -85 405 -65 475
rect -35 405 -15 475
rect -85 150 -65 220
rect -35 150 -15 220
<< metal1 >>
rect -120 575 85 585
rect -120 505 -85 575
rect -65 505 -35 575
rect -15 505 85 575
rect -120 475 85 505
rect -120 405 -85 475
rect -65 405 -35 475
rect -15 405 85 475
rect -120 395 85 405
rect -120 220 85 330
rect -120 150 -85 220
rect -65 150 -35 220
rect -15 150 85 220
rect -120 140 85 150
<< labels >>
rlabel metal1 -120 235 -120 235 7 VN
port 4 w
rlabel locali -25 100 -25 100 7 A
port 1 w
rlabel locali 60 90 60 90 3 Y
port 2 e
rlabel metal1 -120 490 -120 490 7 VP
port 3 w
<< end >>
