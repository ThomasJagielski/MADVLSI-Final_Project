magic
tech sky130A
timestamp 1620437679
<< nwell >>
rect 205 470 415 490
rect 135 250 415 470
<< nmos >>
rect 265 15 280 115
rect 330 15 345 115
<< pmos >>
rect 265 365 280 465
rect 330 365 345 465
<< ndiff >>
rect 215 100 265 115
rect 215 30 230 100
rect 250 30 265 100
rect 215 15 265 30
rect 280 100 330 115
rect 280 30 295 100
rect 315 30 330 100
rect 280 15 330 30
rect 345 100 395 115
rect 345 30 360 100
rect 380 30 395 100
rect 345 15 395 30
<< pdiff >>
rect 215 450 265 465
rect 215 380 230 450
rect 250 380 265 450
rect 215 365 265 380
rect 280 450 330 465
rect 280 380 295 450
rect 315 380 330 450
rect 280 365 330 380
rect 345 450 395 465
rect 345 380 360 450
rect 380 380 395 450
rect 345 365 395 380
<< ndiffc >>
rect 230 30 250 100
rect 295 30 315 100
rect 360 30 380 100
<< pdiffc >>
rect 230 380 250 450
rect 295 380 315 450
rect 360 380 380 450
<< poly >>
rect 95 515 345 525
rect 95 495 105 515
rect 125 510 345 515
rect 125 495 135 510
rect 95 485 135 495
rect 265 465 280 480
rect 330 465 345 510
rect 265 230 280 365
rect 330 350 345 365
rect 160 220 345 230
rect 160 200 170 220
rect 190 215 345 220
rect 190 200 200 215
rect 160 190 200 200
rect 120 125 280 140
rect 265 115 280 125
rect 330 115 345 215
rect 265 0 280 15
rect 330 0 345 15
<< polycont >>
rect 105 495 125 515
rect 170 200 190 220
<< locali >>
rect 0 515 135 525
rect 0 505 105 515
rect 95 495 105 505
rect 125 495 135 515
rect 95 485 135 495
rect 305 505 415 525
rect 305 460 325 505
rect 220 450 260 460
rect 220 380 230 450
rect 250 380 260 450
rect 220 370 260 380
rect 285 450 325 460
rect 285 380 295 450
rect 315 380 325 450
rect 285 370 325 380
rect 350 450 390 460
rect 350 380 360 450
rect 380 380 390 450
rect 350 370 390 380
rect 160 220 200 230
rect 160 200 170 220
rect 190 200 200 220
rect 160 190 200 200
rect 220 110 240 370
rect 285 110 305 370
rect 350 110 370 370
rect 220 100 260 110
rect 220 30 230 100
rect 250 30 260 100
rect 220 20 260 30
rect 285 100 325 110
rect 285 30 295 100
rect 315 30 325 100
rect 285 20 325 30
rect 350 100 390 110
rect 350 30 360 100
rect 380 30 390 100
rect 350 20 390 30
rect 220 -60 240 20
rect 0 -80 240 -60
rect 350 -100 370 20
rect 0 -120 370 -100
<< metal1 >>
rect 205 275 415 465
rect 205 20 415 210
use inverter  inverter_0
timestamp 1620435323
transform 1 0 120 0 1 -120
box -120 80 85 610
<< labels >>
rlabel locali 0 -70 0 -70 7 A
rlabel locali 0 -110 0 -110 7 B
rlabel locali 415 515 415 515 3 muxout
<< end >>
