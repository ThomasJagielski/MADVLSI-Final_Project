magic
tech sky130A
timestamp 1620518861
<< error_p >>
rect 420 4500 480 4650
rect 540 4500 600 4650
rect 660 4500 720 4650
rect 780 4500 840 4650
rect 900 4500 960 4650
rect 1020 4500 1080 4650
rect 1140 4500 1200 4650
rect 1260 4500 1320 4650
rect 1380 4500 1440 4650
rect 420 3300 480 3450
rect 540 3300 600 3450
rect 660 3300 720 3450
rect 780 3300 840 3450
rect 900 3300 960 3450
rect 1020 3300 1080 3450
rect 1140 3300 1200 3450
rect 1260 3300 1320 3450
rect 1380 3300 1440 3450
rect 300 2425 360 2575
rect 420 2425 480 2575
rect 540 2425 600 2575
rect 660 2425 720 2575
rect 780 2425 840 2575
rect 900 2425 960 2575
rect 1020 2425 1080 2575
rect 1140 2425 1200 2575
rect 1260 2425 1320 2575
rect 1380 2425 1440 2575
rect 1500 2425 1560 2575
rect 300 1390 360 1540
rect 420 1390 480 1540
rect 540 1390 600 1540
rect 660 1390 720 1540
rect 780 1390 840 1540
rect 900 1390 960 1540
rect 1020 1390 1080 1540
rect 1140 1390 1200 1540
rect 1260 1390 1320 1540
rect 1380 1390 1440 1540
rect 1500 1390 1560 1540
rect 65 710 115 722
rect 305 710 355 722
rect 545 710 595 722
rect 1265 710 1315 722
rect 1505 710 1555 722
rect 1745 710 1795 722
rect -60 560 0 710
rect 60 560 120 710
rect 180 560 240 710
rect 300 560 360 710
rect 420 560 480 710
rect 540 560 600 710
rect 660 560 720 710
rect 780 560 840 710
rect 900 560 960 710
rect 1020 560 1080 710
rect 1140 560 1200 710
rect 1260 560 1320 710
rect 1380 560 1440 710
rect 1500 560 1560 710
rect 1620 560 1680 710
rect 1740 560 1800 710
rect 1860 560 1920 710
rect -60 0 0 150
rect 60 0 120 150
rect 180 0 240 150
rect 300 0 360 150
rect 420 0 480 150
rect 540 0 600 150
rect 660 0 720 150
rect 780 0 840 150
rect 900 0 960 150
rect 1020 0 1080 150
rect 1140 0 1200 150
rect 1260 0 1320 150
rect 1380 0 1440 150
rect 1500 0 1560 150
rect 1620 0 1680 150
rect 1740 0 1800 150
rect 1860 0 1920 150
<< nmos >>
rect 480 4500 540 4650
rect 600 4500 660 4650
rect 720 4500 780 4650
rect 840 4500 900 4650
rect 960 4500 1020 4650
rect 1080 4500 1140 4650
rect 1200 4500 1260 4650
rect 1320 4500 1380 4650
rect 480 3300 540 3450
rect 600 3300 660 3450
rect 720 3300 780 3450
rect 840 3300 900 3450
rect 960 3300 1020 3450
rect 1080 3300 1140 3450
rect 1200 3300 1260 3450
rect 1320 3300 1380 3450
rect 360 2425 420 2575
rect 480 2425 540 2575
rect 600 2425 660 2575
rect 720 2425 780 2575
rect 840 2425 900 2575
rect 960 2425 1020 2575
rect 1080 2425 1140 2575
rect 1200 2425 1260 2575
rect 1320 2425 1380 2575
rect 1440 2425 1500 2575
rect 360 1390 420 1540
rect 480 1390 540 1540
rect 600 1390 660 1540
rect 720 1390 780 1540
rect 840 1390 900 1540
rect 960 1390 1020 1540
rect 1080 1390 1140 1540
rect 1200 1390 1260 1540
rect 1320 1390 1380 1540
rect 1440 1390 1500 1540
rect 0 560 60 710
rect 120 560 180 710
rect 240 560 300 710
rect 360 560 420 710
rect 480 560 540 710
rect 600 560 660 710
rect 720 560 780 710
rect 840 560 900 710
rect 960 560 1020 710
rect 1080 560 1140 710
rect 1200 560 1260 710
rect 1320 560 1380 710
rect 1440 560 1500 710
rect 1560 560 1620 710
rect 1680 560 1740 710
rect 1800 560 1860 710
rect 0 0 60 150
rect 120 0 180 150
rect 240 0 300 150
rect 360 0 420 150
rect 480 0 540 150
rect 600 0 660 150
rect 720 0 780 150
rect 840 0 900 150
rect 960 0 1020 150
rect 1080 0 1140 150
rect 1200 0 1260 150
rect 1320 0 1380 150
rect 1440 0 1500 150
rect 1560 0 1620 150
rect 1680 0 1740 150
rect 1800 0 1860 150
<< ndiff >>
rect 420 4635 480 4650
rect 420 4515 435 4635
rect 465 4515 480 4635
rect 420 4500 480 4515
rect 540 4635 600 4650
rect 540 4515 555 4635
rect 585 4515 600 4635
rect 540 4500 600 4515
rect 660 4635 720 4650
rect 660 4515 675 4635
rect 705 4515 720 4635
rect 660 4500 720 4515
rect 780 4635 840 4650
rect 780 4515 795 4635
rect 825 4515 840 4635
rect 780 4500 840 4515
rect 900 4635 960 4650
rect 900 4515 915 4635
rect 945 4515 960 4635
rect 900 4500 960 4515
rect 1020 4635 1080 4650
rect 1020 4515 1035 4635
rect 1065 4515 1080 4635
rect 1020 4500 1080 4515
rect 1140 4635 1200 4650
rect 1140 4515 1155 4635
rect 1185 4515 1200 4635
rect 1140 4500 1200 4515
rect 1260 4635 1320 4650
rect 1260 4515 1275 4635
rect 1305 4515 1320 4635
rect 1260 4500 1320 4515
rect 1380 4635 1440 4650
rect 1380 4515 1395 4635
rect 1425 4515 1440 4635
rect 1380 4500 1440 4515
rect 420 3435 480 3450
rect 420 3315 435 3435
rect 465 3315 480 3435
rect 420 3300 480 3315
rect 540 3435 600 3450
rect 540 3315 555 3435
rect 585 3315 600 3435
rect 540 3300 600 3315
rect 660 3435 720 3450
rect 660 3315 675 3435
rect 705 3315 720 3435
rect 660 3300 720 3315
rect 780 3435 840 3450
rect 780 3315 795 3435
rect 825 3315 840 3435
rect 780 3300 840 3315
rect 900 3435 960 3450
rect 900 3315 915 3435
rect 945 3315 960 3435
rect 900 3300 960 3315
rect 1020 3435 1080 3450
rect 1020 3315 1035 3435
rect 1065 3315 1080 3435
rect 1020 3300 1080 3315
rect 1140 3435 1200 3450
rect 1140 3315 1155 3435
rect 1185 3315 1200 3435
rect 1140 3300 1200 3315
rect 1260 3435 1320 3450
rect 1260 3315 1275 3435
rect 1305 3315 1320 3435
rect 1260 3300 1320 3315
rect 1380 3435 1440 3450
rect 1380 3315 1395 3435
rect 1425 3315 1440 3435
rect 1380 3300 1440 3315
rect 300 2560 360 2575
rect 300 2440 315 2560
rect 345 2440 360 2560
rect 300 2425 360 2440
rect 420 2560 480 2575
rect 420 2440 435 2560
rect 465 2440 480 2560
rect 420 2425 480 2440
rect 540 2560 600 2575
rect 540 2440 555 2560
rect 585 2440 600 2560
rect 540 2425 600 2440
rect 660 2560 720 2575
rect 660 2440 675 2560
rect 705 2440 720 2560
rect 660 2425 720 2440
rect 780 2560 840 2575
rect 780 2440 795 2560
rect 825 2440 840 2560
rect 780 2425 840 2440
rect 900 2560 960 2575
rect 900 2440 915 2560
rect 945 2440 960 2560
rect 900 2425 960 2440
rect 1020 2560 1080 2575
rect 1020 2440 1035 2560
rect 1065 2440 1080 2560
rect 1020 2425 1080 2440
rect 1140 2560 1200 2575
rect 1140 2440 1155 2560
rect 1185 2440 1200 2560
rect 1140 2425 1200 2440
rect 1260 2560 1320 2575
rect 1260 2440 1275 2560
rect 1305 2440 1320 2560
rect 1260 2425 1320 2440
rect 1380 2560 1440 2575
rect 1380 2440 1395 2560
rect 1425 2440 1440 2560
rect 1380 2425 1440 2440
rect 1500 2560 1560 2575
rect 1500 2440 1515 2560
rect 1545 2440 1560 2560
rect 1500 2425 1560 2440
rect 300 1525 360 1540
rect 300 1405 315 1525
rect 345 1405 360 1525
rect 300 1390 360 1405
rect 420 1525 480 1540
rect 420 1405 435 1525
rect 465 1405 480 1525
rect 420 1390 480 1405
rect 540 1525 600 1540
rect 540 1405 555 1525
rect 585 1405 600 1525
rect 540 1390 600 1405
rect 660 1525 720 1540
rect 660 1405 675 1525
rect 705 1405 720 1525
rect 660 1390 720 1405
rect 780 1525 840 1540
rect 780 1405 795 1525
rect 825 1405 840 1525
rect 780 1390 840 1405
rect 900 1525 960 1540
rect 900 1405 915 1525
rect 945 1405 960 1525
rect 900 1390 960 1405
rect 1020 1525 1080 1540
rect 1020 1405 1035 1525
rect 1065 1405 1080 1525
rect 1020 1390 1080 1405
rect 1140 1525 1200 1540
rect 1140 1405 1155 1525
rect 1185 1405 1200 1525
rect 1140 1390 1200 1405
rect 1260 1525 1320 1540
rect 1260 1405 1275 1525
rect 1305 1405 1320 1525
rect 1260 1390 1320 1405
rect 1380 1525 1440 1540
rect 1380 1405 1395 1525
rect 1425 1405 1440 1525
rect 1380 1390 1440 1405
rect 1500 1525 1560 1540
rect 1500 1405 1515 1525
rect 1545 1405 1560 1525
rect 1500 1390 1560 1405
rect -60 695 0 710
rect -60 575 -45 695
rect -15 575 0 695
rect -60 560 0 575
rect 60 695 120 710
rect 60 575 75 695
rect 105 575 120 695
rect 60 560 120 575
rect 180 695 240 710
rect 180 575 195 695
rect 225 575 240 695
rect 180 560 240 575
rect 300 695 360 710
rect 300 575 315 695
rect 345 575 360 695
rect 300 560 360 575
rect 420 695 480 710
rect 420 575 435 695
rect 465 575 480 695
rect 420 560 480 575
rect 540 695 600 710
rect 540 575 555 695
rect 585 575 600 695
rect 540 560 600 575
rect 660 695 720 710
rect 660 575 675 695
rect 705 575 720 695
rect 660 560 720 575
rect 780 695 840 710
rect 780 575 795 695
rect 825 575 840 695
rect 780 560 840 575
rect 900 695 960 710
rect 900 575 915 695
rect 945 575 960 695
rect 900 560 960 575
rect 1020 695 1080 710
rect 1020 575 1035 695
rect 1065 575 1080 695
rect 1020 560 1080 575
rect 1140 695 1200 710
rect 1140 575 1155 695
rect 1185 575 1200 695
rect 1140 560 1200 575
rect 1260 695 1320 710
rect 1260 575 1275 695
rect 1305 575 1320 695
rect 1260 560 1320 575
rect 1380 695 1440 710
rect 1380 575 1395 695
rect 1425 575 1440 695
rect 1380 560 1440 575
rect 1500 695 1560 710
rect 1500 575 1515 695
rect 1545 575 1560 695
rect 1500 560 1560 575
rect 1620 695 1680 710
rect 1620 575 1635 695
rect 1665 575 1680 695
rect 1620 560 1680 575
rect 1740 695 1800 710
rect 1740 575 1755 695
rect 1785 575 1800 695
rect 1740 560 1800 575
rect 1860 695 1920 710
rect 1860 575 1875 695
rect 1905 575 1920 695
rect 1860 560 1920 575
rect -60 135 0 150
rect -60 15 -45 135
rect -15 15 0 135
rect -60 0 0 15
rect 60 135 120 150
rect 60 15 75 135
rect 105 15 120 135
rect 60 0 120 15
rect 180 135 240 150
rect 180 15 195 135
rect 225 15 240 135
rect 180 0 240 15
rect 300 135 360 150
rect 300 15 315 135
rect 345 15 360 135
rect 300 0 360 15
rect 420 135 480 150
rect 420 15 435 135
rect 465 15 480 135
rect 420 0 480 15
rect 540 135 600 150
rect 540 15 555 135
rect 585 15 600 135
rect 540 0 600 15
rect 660 135 720 150
rect 660 15 675 135
rect 705 15 720 135
rect 660 0 720 15
rect 780 135 840 150
rect 780 15 795 135
rect 825 15 840 135
rect 780 0 840 15
rect 900 135 960 150
rect 900 15 915 135
rect 945 15 960 135
rect 900 0 960 15
rect 1020 135 1080 150
rect 1020 15 1035 135
rect 1065 15 1080 135
rect 1020 0 1080 15
rect 1140 135 1200 150
rect 1140 15 1155 135
rect 1185 15 1200 135
rect 1140 0 1200 15
rect 1260 135 1320 150
rect 1260 15 1275 135
rect 1305 15 1320 135
rect 1260 0 1320 15
rect 1380 135 1440 150
rect 1380 15 1395 135
rect 1425 15 1440 135
rect 1380 0 1440 15
rect 1500 135 1560 150
rect 1500 15 1515 135
rect 1545 15 1560 135
rect 1500 0 1560 15
rect 1620 135 1680 150
rect 1620 15 1635 135
rect 1665 15 1680 135
rect 1620 0 1680 15
rect 1740 135 1800 150
rect 1740 15 1755 135
rect 1785 15 1800 135
rect 1740 0 1800 15
rect 1860 135 1920 150
rect 1860 15 1875 135
rect 1905 15 1920 135
rect 1860 0 1920 15
<< ndiffc >>
rect 435 4515 465 4635
rect 555 4515 585 4635
rect 675 4515 705 4635
rect 795 4515 825 4635
rect 915 4515 945 4635
rect 1035 4515 1065 4635
rect 1155 4515 1185 4635
rect 1275 4515 1305 4635
rect 1395 4515 1425 4635
rect 435 3315 465 3435
rect 555 3315 585 3435
rect 675 3315 705 3435
rect 795 3315 825 3435
rect 915 3315 945 3435
rect 1035 3315 1065 3435
rect 1155 3315 1185 3435
rect 1275 3315 1305 3435
rect 1395 3315 1425 3435
rect 315 2440 345 2560
rect 435 2440 465 2560
rect 555 2440 585 2560
rect 675 2440 705 2560
rect 795 2440 825 2560
rect 915 2440 945 2560
rect 1035 2440 1065 2560
rect 1155 2440 1185 2560
rect 1275 2440 1305 2560
rect 1395 2440 1425 2560
rect 1515 2440 1545 2560
rect 315 1405 345 1525
rect 435 1405 465 1525
rect 555 1405 585 1525
rect 675 1405 705 1525
rect 795 1405 825 1525
rect 915 1405 945 1525
rect 1035 1405 1065 1525
rect 1155 1405 1185 1525
rect 1275 1405 1305 1525
rect 1395 1405 1425 1525
rect 1515 1405 1545 1525
rect -45 575 -15 695
rect 75 575 105 695
rect 195 575 225 695
rect 315 575 345 695
rect 435 575 465 695
rect 555 575 585 695
rect 675 575 705 695
rect 795 575 825 695
rect 915 575 945 695
rect 1035 575 1065 695
rect 1155 575 1185 695
rect 1275 575 1305 695
rect 1395 575 1425 695
rect 1515 575 1545 695
rect 1635 575 1665 695
rect 1755 575 1785 695
rect 1875 575 1905 695
rect -45 15 -15 135
rect 75 15 105 135
rect 195 15 225 135
rect 315 15 345 135
rect 435 15 465 135
rect 555 15 585 135
rect 675 15 705 135
rect 795 15 825 135
rect 915 15 945 135
rect 1035 15 1065 135
rect 1155 15 1185 135
rect 1275 15 1305 135
rect 1395 15 1425 135
rect 1515 15 1545 135
rect 1635 15 1665 135
rect 1755 15 1785 135
rect 1875 15 1905 135
<< poly >>
rect 420 4690 1380 4705
rect 480 4650 540 4690
rect 600 4650 660 4665
rect 720 4650 780 4665
rect 840 4650 900 4665
rect 960 4650 1020 4665
rect 1080 4650 1140 4665
rect 1200 4650 1260 4665
rect 1320 4650 1380 4690
rect 480 3450 540 4500
rect 600 4485 660 4500
rect 720 4460 780 4500
rect 600 4445 780 4460
rect 600 3450 660 4445
rect 840 4420 900 4500
rect 960 4420 1020 4500
rect 1080 4460 1140 4500
rect 1200 4485 1260 4500
rect 1080 4445 1260 4460
rect 840 4405 1020 4420
rect 720 3450 780 3465
rect 840 3450 900 3465
rect 960 3450 1020 3465
rect 1080 3450 1140 3465
rect 1200 3450 1260 4445
rect 1320 3450 1380 4500
rect 480 3285 540 3300
rect 600 3260 660 3300
rect 720 3285 780 3300
rect 420 3245 660 3260
rect 840 3260 900 3300
rect 960 3260 1020 3300
rect 1080 3285 1140 3300
rect 1200 3285 1260 3300
rect 1320 3285 1380 3300
rect 840 3245 1020 3260
rect 360 2615 1500 2630
rect 360 2575 420 2615
rect 480 2575 540 2590
rect 600 2575 660 2590
rect 720 2575 780 2615
rect 840 2575 900 2590
rect 960 2575 1020 2590
rect 1080 2575 1140 2615
rect 1200 2575 1260 2590
rect 1320 2575 1380 2590
rect 1440 2575 1500 2615
rect 360 2410 420 2425
rect 480 2400 540 2425
rect 600 2410 660 2425
rect 720 2410 780 2425
rect 480 2380 490 2400
rect 530 2380 540 2400
rect 480 2370 540 2380
rect 840 2400 900 2425
rect 840 2380 850 2400
rect 890 2380 900 2400
rect 840 2370 900 2380
rect 960 2400 1020 2425
rect 1080 2410 1140 2425
rect 1200 2410 1260 2425
rect 960 2380 970 2400
rect 1010 2380 1020 2400
rect 960 2370 1020 2380
rect 1320 2400 1380 2425
rect 1440 2410 1500 2425
rect 1320 2380 1330 2400
rect 1370 2380 1380 2400
rect 1320 2370 1380 2380
rect 910 2340 950 2350
rect 910 2320 920 2340
rect 940 2320 950 2340
rect 910 2310 950 2320
rect 920 1655 940 2310
rect 910 1645 950 1655
rect 910 1625 920 1645
rect 940 1625 950 1645
rect 910 1615 950 1625
rect 480 1585 540 1595
rect 480 1565 490 1585
rect 530 1565 540 1585
rect 360 1540 420 1555
rect 480 1540 540 1565
rect 840 1585 900 1595
rect 840 1565 850 1585
rect 890 1565 900 1585
rect 600 1540 660 1555
rect 720 1540 780 1555
rect 840 1540 900 1565
rect 960 1585 1020 1595
rect 960 1565 970 1585
rect 1010 1565 1020 1585
rect 960 1540 1020 1565
rect 1320 1585 1380 1595
rect 1320 1565 1330 1585
rect 1370 1565 1380 1585
rect 1080 1540 1140 1555
rect 1200 1540 1260 1555
rect 1320 1540 1380 1565
rect 1440 1540 1500 1555
rect 360 1350 420 1390
rect 480 1375 540 1390
rect 600 1375 660 1390
rect 720 1350 780 1390
rect 840 1375 900 1390
rect 960 1375 1020 1390
rect 1080 1350 1140 1390
rect 1200 1375 1260 1390
rect 1320 1375 1380 1390
rect 1440 1350 1500 1390
rect 360 1335 1500 1350
rect 0 710 60 725
rect 120 710 180 725
rect 240 710 300 725
rect 360 710 420 725
rect 480 710 540 725
rect 600 710 660 725
rect 720 710 780 725
rect 840 710 900 725
rect 960 710 1020 725
rect 1080 710 1140 725
rect 1200 710 1260 725
rect 1320 710 1380 725
rect 1440 710 1500 725
rect 1560 710 1620 725
rect 1680 710 1740 725
rect 1800 710 1860 725
rect 0 520 60 560
rect 120 520 180 560
rect 240 520 300 560
rect 360 545 420 560
rect 480 520 540 560
rect 600 520 660 560
rect 720 545 780 560
rect 840 520 900 560
rect 960 520 1020 560
rect 1080 545 1140 560
rect 1200 520 1260 560
rect 1320 520 1380 560
rect 1440 545 1500 560
rect 1560 520 1620 560
rect 1680 520 1740 560
rect 1800 520 1860 560
rect 0 505 1860 520
rect 785 470 835 480
rect 785 445 795 470
rect 825 450 835 470
rect 1030 470 1080 480
rect 1030 450 1040 470
rect 825 445 1040 450
rect 1070 445 1080 470
rect 425 430 475 445
rect 785 435 1080 445
rect 425 405 435 430
rect 465 410 475 430
rect 1385 430 1435 445
rect 1385 410 1395 430
rect 465 405 1395 410
rect 1425 405 1435 430
rect 425 395 1435 405
rect 0 150 60 165
rect 120 150 180 165
rect 240 150 300 165
rect 360 150 420 165
rect 480 150 540 165
rect 600 150 660 165
rect 720 150 780 165
rect 840 150 900 165
rect 960 150 1020 165
rect 1080 150 1140 165
rect 1200 150 1260 165
rect 1320 150 1380 165
rect 1440 150 1500 165
rect 1560 150 1620 165
rect 1680 150 1740 165
rect 1800 150 1860 165
rect 0 -40 60 0
rect 120 -40 180 0
rect 240 -40 300 0
rect 360 -15 420 0
rect 480 -40 540 0
rect 600 -40 660 0
rect 720 -15 780 0
rect 840 -40 900 0
rect 960 -40 1020 0
rect 1080 -15 1140 0
rect 1200 -40 1260 0
rect 1320 -40 1380 0
rect 1440 -15 1500 0
rect 1560 -40 1620 0
rect 1680 -40 1740 0
rect 1800 -40 1860 0
rect 0 -55 1860 -40
<< polycont >>
rect 490 2380 530 2400
rect 850 2380 890 2400
rect 970 2380 1010 2400
rect 1330 2380 1370 2400
rect 920 2320 940 2340
rect 920 1625 940 1645
rect 490 1565 530 1585
rect 850 1565 890 1585
rect 970 1565 1010 1585
rect 1330 1565 1370 1585
rect 795 445 825 470
rect 1040 445 1070 470
rect 435 405 465 430
rect 1395 405 1425 430
<< locali >>
rect 425 4850 1435 4870
rect 425 4635 475 4850
rect 425 4515 435 4635
rect 465 4515 475 4635
rect 425 4505 475 4515
rect 545 4810 1315 4830
rect 545 4635 595 4810
rect 545 4515 555 4635
rect 585 4515 595 4635
rect 545 4505 595 4515
rect 665 4635 715 4645
rect 665 4515 675 4635
rect 705 4515 715 4635
rect 665 4320 715 4515
rect 785 4635 835 4810
rect 785 4515 795 4635
rect 825 4515 835 4635
rect 785 4505 835 4515
rect 905 4635 955 4645
rect 905 4515 915 4635
rect 945 4515 955 4635
rect 905 4505 955 4515
rect 1025 4635 1075 4810
rect 1025 4515 1035 4635
rect 1065 4515 1075 4635
rect 1025 4505 1075 4515
rect 1145 4635 1195 4645
rect 1145 4515 1155 4635
rect 1185 4515 1195 4635
rect 1145 4320 1195 4515
rect 1265 4635 1315 4810
rect 1265 4515 1275 4635
rect 1305 4515 1315 4635
rect 1265 4505 1315 4515
rect 1385 4635 1435 4850
rect 1385 4515 1395 4635
rect 1425 4515 1435 4635
rect 1385 4505 1435 4515
rect 665 4300 1195 4320
rect 665 3635 1195 3655
rect 425 3435 475 3445
rect 425 3315 435 3435
rect 465 3315 475 3435
rect 425 3095 475 3315
rect 545 3435 595 3445
rect 545 3315 555 3435
rect 585 3315 595 3435
rect 545 3135 595 3315
rect 665 3435 715 3635
rect 665 3315 675 3435
rect 705 3315 715 3435
rect 665 3305 715 3315
rect 785 3435 835 3445
rect 785 3315 795 3435
rect 825 3315 835 3435
rect 785 3135 835 3315
rect 905 3435 955 3445
rect 905 3315 915 3435
rect 945 3315 955 3435
rect 905 3305 955 3315
rect 1025 3435 1075 3445
rect 1025 3315 1035 3435
rect 1065 3315 1075 3435
rect 1025 3135 1075 3315
rect 1145 3435 1195 3635
rect 1145 3315 1155 3435
rect 1185 3315 1195 3435
rect 1145 3305 1195 3315
rect 1265 3435 1315 3445
rect 1265 3315 1275 3435
rect 1305 3315 1315 3435
rect 1265 3135 1315 3315
rect 545 3115 1315 3135
rect 1385 3435 1435 3445
rect 1385 3315 1395 3435
rect 1425 3315 1435 3435
rect 1385 3095 1435 3315
rect 425 3075 1435 3095
rect 425 2840 1435 2860
rect 305 2560 355 2570
rect 305 2440 315 2560
rect 345 2440 355 2560
rect 305 2430 355 2440
rect 425 2560 475 2840
rect 785 2660 1075 2680
rect 425 2440 435 2560
rect 465 2440 475 2560
rect 425 2430 475 2440
rect 545 2560 595 2570
rect 545 2440 555 2560
rect 585 2440 595 2560
rect 545 2410 595 2440
rect 665 2560 715 2570
rect 665 2440 675 2560
rect 705 2440 715 2560
rect 665 2430 715 2440
rect 785 2560 835 2660
rect 785 2440 795 2560
rect 825 2440 835 2560
rect 785 2430 835 2440
rect 905 2560 955 2570
rect 905 2440 915 2560
rect 945 2440 955 2560
rect 905 2430 955 2440
rect 1025 2560 1075 2660
rect 1025 2440 1035 2560
rect 1065 2440 1075 2560
rect 1025 2430 1075 2440
rect 1145 2560 1195 2570
rect 1145 2440 1155 2560
rect 1185 2440 1195 2560
rect 1145 2430 1195 2440
rect 1265 2560 1315 2570
rect 1265 2440 1275 2560
rect 1305 2440 1315 2560
rect 480 2400 595 2410
rect 480 2380 490 2400
rect 530 2380 595 2400
rect 480 2370 595 2380
rect 840 2400 900 2410
rect 840 2380 850 2400
rect 890 2380 900 2400
rect 840 2370 900 2380
rect 480 2205 540 2370
rect 840 2205 890 2370
rect 920 2350 940 2430
rect 1265 2410 1315 2440
rect 1385 2560 1435 2840
rect 1385 2440 1395 2560
rect 1425 2440 1435 2560
rect 1385 2430 1435 2440
rect 1505 2560 1555 2570
rect 1505 2440 1515 2560
rect 1545 2440 1555 2560
rect 1505 2430 1555 2440
rect 960 2400 1020 2410
rect 960 2380 970 2400
rect 1010 2380 1020 2400
rect 960 2370 1020 2380
rect 1265 2400 1380 2410
rect 1265 2380 1330 2400
rect 1370 2380 1380 2400
rect 1265 2370 1380 2380
rect 910 2340 950 2350
rect 910 2320 920 2340
rect 940 2320 950 2340
rect 910 2310 950 2320
rect 970 2205 1020 2370
rect 1320 2205 1380 2370
rect 480 2185 1380 2205
rect 480 1595 540 2185
rect 840 1595 890 2185
rect 910 1645 950 1655
rect 910 1625 920 1645
rect 940 1625 950 1645
rect 910 1615 950 1625
rect 480 1585 595 1595
rect 480 1565 490 1585
rect 530 1565 595 1585
rect 480 1555 595 1565
rect 840 1585 900 1595
rect 840 1565 850 1585
rect 890 1565 900 1585
rect 840 1555 900 1565
rect 305 1525 355 1535
rect 305 1405 315 1525
rect 345 1405 355 1525
rect 305 1395 355 1405
rect 425 1525 475 1535
rect 425 1405 435 1525
rect 465 1405 475 1525
rect 425 1120 475 1405
rect 545 1525 595 1555
rect 920 1535 940 1615
rect 970 1595 1020 2185
rect 1320 1595 1380 2185
rect 960 1585 1020 1595
rect 960 1565 970 1585
rect 1010 1565 1020 1585
rect 960 1555 1020 1565
rect 1265 1585 1380 1595
rect 1265 1565 1330 1585
rect 1370 1565 1380 1585
rect 1265 1555 1380 1565
rect 545 1405 555 1525
rect 585 1405 595 1525
rect 545 1395 595 1405
rect 665 1525 715 1535
rect 665 1405 675 1525
rect 705 1405 715 1525
rect 665 1395 715 1405
rect 785 1525 835 1535
rect 785 1405 795 1525
rect 825 1405 835 1525
rect 785 1300 835 1405
rect 905 1525 955 1535
rect 905 1405 915 1525
rect 945 1405 955 1525
rect 905 1395 955 1405
rect 1025 1525 1075 1535
rect 1025 1405 1035 1525
rect 1065 1405 1075 1525
rect 1025 1300 1075 1405
rect 1145 1525 1195 1535
rect 1145 1405 1155 1525
rect 1185 1405 1195 1525
rect 1145 1395 1195 1405
rect 1265 1525 1315 1555
rect 1265 1405 1275 1525
rect 1305 1405 1315 1525
rect 1265 1395 1315 1405
rect 1385 1525 1435 1535
rect 1385 1405 1395 1525
rect 1425 1405 1435 1525
rect 785 1280 1075 1300
rect 1385 1120 1435 1405
rect 1505 1525 1555 1535
rect 1505 1405 1515 1525
rect 1545 1405 1555 1525
rect 1505 1395 1555 1405
rect 425 1100 1435 1120
rect 65 805 1795 825
rect 65 710 115 805
rect 305 710 355 805
rect 545 710 595 805
rect 1265 710 1315 805
rect 1505 710 1555 805
rect 1745 710 1795 805
rect -55 695 -5 705
rect -55 575 -45 695
rect -15 575 -5 695
rect -55 565 -5 575
rect 65 695 115 705
rect 65 575 75 695
rect 105 575 115 695
rect 65 565 115 575
rect 185 695 235 705
rect 185 575 195 695
rect 225 575 235 695
rect 185 565 235 575
rect 305 695 355 705
rect 305 575 315 695
rect 345 575 355 695
rect 305 565 355 575
rect 425 695 475 705
rect 425 575 435 695
rect 465 575 475 695
rect 425 430 475 575
rect 545 695 595 705
rect 545 575 555 695
rect 585 575 595 695
rect 545 565 595 575
rect 665 695 715 705
rect 665 575 675 695
rect 705 575 715 695
rect 665 565 715 575
rect 785 695 835 705
rect 785 575 795 695
rect 825 575 835 695
rect 785 470 835 575
rect 785 445 795 470
rect 825 445 835 470
rect 785 435 835 445
rect 905 695 955 705
rect 905 575 915 695
rect 945 575 955 695
rect 425 405 435 430
rect 465 405 475 430
rect 425 395 475 405
rect 905 350 955 575
rect 1025 695 1075 705
rect 1025 575 1035 695
rect 1065 575 1075 695
rect 1025 565 1075 575
rect 1145 695 1195 705
rect 1145 575 1155 695
rect 1185 575 1195 695
rect 1145 565 1195 575
rect 1265 695 1315 705
rect 1265 575 1275 695
rect 1305 575 1315 695
rect 1265 565 1315 575
rect 1385 695 1435 705
rect 1385 575 1395 695
rect 1425 575 1435 695
rect 1030 470 1080 565
rect 1030 445 1040 470
rect 1070 445 1080 470
rect 1030 435 1080 445
rect 1385 430 1435 575
rect 1505 695 1555 705
rect 1505 575 1515 695
rect 1545 575 1555 695
rect 1505 565 1555 575
rect 1625 695 1675 705
rect 1625 575 1635 695
rect 1665 575 1675 695
rect 1625 565 1675 575
rect 1745 695 1795 705
rect 1745 575 1755 695
rect 1785 575 1795 695
rect 1745 565 1795 575
rect 1865 695 1915 705
rect 1865 575 1875 695
rect 1905 575 1915 695
rect 1865 565 1915 575
rect 1385 405 1395 430
rect 1425 405 1435 430
rect 1385 395 1435 405
rect 665 330 1195 350
rect -55 135 -5 145
rect -55 15 -45 135
rect -15 15 -5 135
rect -55 5 -5 15
rect 65 135 115 145
rect 65 15 75 135
rect 105 15 115 135
rect 65 -95 115 15
rect 185 135 235 145
rect 185 15 195 135
rect 225 15 235 135
rect 185 5 235 15
rect 305 135 355 145
rect 305 15 315 135
rect 345 15 355 135
rect 305 -95 355 15
rect 425 135 475 145
rect 425 15 435 135
rect 465 15 475 135
rect 425 5 475 15
rect 545 135 595 145
rect 545 15 555 135
rect 585 15 595 135
rect 545 -95 595 15
rect 665 135 715 330
rect 665 15 675 135
rect 705 15 715 135
rect 665 5 715 15
rect 785 190 1075 210
rect 785 135 835 190
rect 785 15 795 135
rect 825 15 835 135
rect 785 5 835 15
rect 905 135 955 145
rect 905 15 915 135
rect 945 15 955 135
rect 905 5 955 15
rect 1025 135 1075 190
rect 1025 15 1035 135
rect 1065 15 1075 135
rect 1025 5 1075 15
rect 1145 135 1195 330
rect 1145 15 1155 135
rect 1185 15 1195 135
rect 1145 5 1195 15
rect 1265 135 1315 145
rect 1265 15 1275 135
rect 1305 15 1315 135
rect 1265 -95 1315 15
rect 1385 135 1435 145
rect 1385 15 1395 135
rect 1425 15 1435 135
rect 1385 5 1435 15
rect 1505 135 1555 145
rect 1505 15 1515 135
rect 1545 15 1555 135
rect 1505 -95 1555 15
rect 1625 135 1675 145
rect 1625 15 1635 135
rect 1665 15 1675 135
rect 1625 5 1675 15
rect 1745 135 1795 145
rect 1745 15 1755 135
rect 1785 15 1795 135
rect 1745 -95 1795 15
rect 1865 135 1915 145
rect 1865 15 1875 135
rect 1905 15 1915 135
rect 1865 5 1915 15
rect 65 -115 1795 -95
<< end >>
