magic
tech sky130A
timestamp 1620696597
<< nwell >>
rect -110 345 245 590
<< nmos >>
rect -40 75 -25 175
rect 35 75 50 275
rect 110 75 125 175
<< pmos >>
rect -40 470 -25 570
rect 35 370 50 570
rect 110 470 125 570
<< ndiff >>
rect -15 260 35 275
rect -15 175 0 260
rect -90 160 -40 175
rect -90 90 -75 160
rect -55 90 -40 160
rect -90 75 -40 90
rect -25 90 0 175
rect 20 90 35 260
rect -25 75 35 90
rect 50 260 100 275
rect 50 90 65 260
rect 85 175 100 260
rect 85 90 110 175
rect 50 75 110 90
rect 125 160 175 175
rect 125 90 140 160
rect 160 90 175 160
rect 125 75 175 90
<< pdiff >>
rect -90 555 -40 570
rect -90 485 -75 555
rect -55 485 -40 555
rect -90 470 -40 485
rect -25 555 35 570
rect -25 470 0 555
rect -15 385 0 470
rect 20 385 35 555
rect -15 370 35 385
rect 50 555 110 570
rect 50 385 65 555
rect 85 470 110 555
rect 125 555 175 570
rect 125 485 140 555
rect 160 485 175 555
rect 125 470 175 485
rect 85 385 100 470
rect 50 370 100 385
<< ndiffc >>
rect -75 90 -55 160
rect 0 90 20 260
rect 65 90 85 260
rect 140 90 160 160
<< pdiffc >>
rect -75 485 -55 555
rect 0 385 20 555
rect 65 385 85 555
rect 140 485 160 555
<< psubdiff >>
rect 175 160 225 175
rect 175 90 190 160
rect 210 90 225 160
rect 175 75 225 90
<< nsubdiff >>
rect 175 555 225 570
rect 175 485 190 555
rect 210 485 225 555
rect 175 470 225 485
<< psubdiffcont >>
rect 190 90 210 160
<< nsubdiffcont >>
rect 190 485 210 555
<< poly >>
rect -90 615 125 625
rect -90 595 -80 615
rect -60 610 125 615
rect -60 595 -25 610
rect -90 585 -25 595
rect -40 570 -25 585
rect 35 570 50 585
rect 110 570 125 610
rect -40 455 -25 470
rect 35 355 50 370
rect -40 340 50 355
rect -40 175 -25 340
rect 110 330 125 470
rect 70 315 125 330
rect 70 305 85 315
rect 35 290 85 305
rect 35 275 50 290
rect 110 175 125 290
rect -40 60 -25 75
rect 35 60 50 75
rect -90 50 -25 60
rect -90 30 -80 50
rect -60 35 -25 50
rect 110 35 125 75
rect -60 30 125 35
rect -90 20 125 30
<< polycont >>
rect -80 595 -60 615
rect -80 30 -60 50
<< locali >>
rect -90 615 -50 625
rect -90 595 -80 615
rect -60 595 -50 615
rect -90 585 -50 595
rect -85 555 30 565
rect -85 485 -75 555
rect -55 485 0 555
rect -85 475 0 485
rect -10 385 0 475
rect 20 385 30 555
rect -10 340 30 385
rect -110 300 30 340
rect -10 260 30 300
rect -10 170 0 260
rect -85 160 0 170
rect -85 90 -75 160
rect -55 90 0 160
rect 20 90 30 260
rect -85 80 30 90
rect 55 555 220 565
rect 55 385 65 555
rect 85 485 140 555
rect 160 485 190 555
rect 210 485 220 555
rect 85 475 220 485
rect 85 385 95 475
rect 55 340 95 385
rect 55 300 245 340
rect 55 260 95 300
rect 55 90 65 260
rect 85 170 95 260
rect 85 160 220 170
rect 85 90 140 160
rect 160 90 190 160
rect 210 90 220 160
rect 55 80 220 90
rect -90 50 -50 60
rect -90 30 -80 50
rect -60 30 -50 50
rect -90 20 -50 30
<< labels >>
rlabel locali -90 40 -90 40 7 nCLK
rlabel locali -90 605 -90 605 7 CLK
rlabel locali 245 320 245 320 3 B
rlabel locali -110 320 -110 320 7 A
<< end >>
