magic
tech sky130A
timestamp 1620771670
<< poly >>
rect -160 10875 210 10885
rect -160 10855 -150 10875
rect -130 10870 180 10875
rect -130 10855 -120 10870
rect -160 10845 -120 10855
rect 170 10855 180 10870
rect 200 10855 210 10875
rect 170 10845 210 10855
rect -115 8715 -70 8725
rect -115 8695 -105 8715
rect -80 8695 -70 8715
rect -115 8685 -70 8695
rect 33410 5715 33510 5725
rect 33410 5695 33420 5715
rect 33440 5710 33510 5715
rect 33440 5695 33450 5710
rect 33410 5685 33450 5695
<< polycont >>
rect -150 10855 -130 10875
rect 180 10855 200 10875
rect -105 8695 -80 8715
rect 33420 5695 33440 5715
<< locali >>
rect -140 18005 10010 18025
rect -140 10885 -120 18005
rect -160 10875 -120 10885
rect -160 10855 -150 10875
rect -130 10855 -120 10875
rect -160 10845 -120 10855
rect -100 17965 5045 17985
rect -100 8725 -80 17965
rect 5025 17920 5045 17965
rect -60 17255 15 17275
rect -60 10985 -40 17255
rect -60 10945 155 10985
rect 170 10875 210 10885
rect 170 10855 180 10875
rect 200 10855 210 10875
rect 170 10845 210 10855
rect -115 8715 -70 8725
rect -115 8695 -105 8715
rect -80 8695 -70 8715
rect -115 8685 -70 8695
rect 27555 5745 33495 5765
rect 27555 5725 27690 5745
rect 27555 5705 27575 5725
rect 27970 5715 33450 5725
rect 27970 5705 33420 5715
rect 33410 5695 33420 5705
rect 33440 5695 33450 5715
rect 33410 5685 33450 5695
rect 27470 5120 27585 5140
rect 27470 5080 27500 5120
rect 32120 -2475 32160 -2420
rect 33475 -2475 33495 5745
rect 32120 -2495 33495 -2475
<< viali >>
rect -105 8695 -80 8715
rect 27915 5280 27935 5300
<< metal1 >>
rect 10350 11720 31365 11805
rect 7185 11610 31365 11720
rect 7185 11015 23110 11610
rect 7185 10965 18775 11015
rect -115 8720 -70 8725
rect -115 8690 -110 8720
rect -75 8690 -70 8720
rect -115 8685 -70 8690
rect 27970 5650 28175 5665
rect 27970 5490 27985 5650
rect 28160 5490 28175 5650
rect 27970 5475 28175 5490
rect 30995 5410 31365 11610
rect 27970 5220 31365 5410
rect 30995 4515 31365 5220
rect 30965 3980 31365 4515
rect 30995 15 31365 3980
rect 30995 -520 34065 15
rect 33425 -1080 33525 -1075
rect 33425 -1260 33480 -1080
rect 33520 -1260 33525 -1080
rect 33425 -1265 33525 -1260
rect 33695 -1330 34065 -520
rect 33255 -1520 34065 -1330
rect 33705 -1990 34065 -1520
rect 33455 -2180 34065 -1990
<< via1 >>
rect -110 8715 -75 8720
rect -110 8695 -105 8715
rect -105 8695 -80 8715
rect -80 8695 -75 8715
rect -110 8690 -75 8695
rect 27985 5490 28160 5650
rect 33480 -1260 33520 -1080
<< metal2 >>
rect 10265 11890 31365 12080
rect -115 8720 -70 8725
rect -115 8690 -110 8720
rect -75 8690 -70 8720
rect -115 8685 -70 8690
rect 27975 5650 28170 5660
rect 27975 5490 27985 5650
rect 28160 5490 28170 5650
rect 27975 4525 28170 5490
rect 30995 4525 31365 11890
rect 22650 3975 31365 4525
rect 30995 15 31365 3975
rect 30995 -520 34065 15
rect 33695 -1075 34065 -520
rect 33475 -1080 34065 -1075
rect 33475 -1260 33480 -1080
rect 33520 -1260 34065 -1080
rect 33475 -1265 34065 -1260
<< via2 >>
rect -110 8690 -75 8720
<< metal3 >>
rect -120 8720 5 8735
rect -120 8690 -110 8720
rect -75 8690 5 8720
rect -120 8680 5 8690
use adc  adc_0
timestamp 1620769246
transform 1 0 8045 0 1 -4180
box -7870 -175 25410 3310
use mux2  mux2_0
timestamp 1620437679
transform 1 0 27555 0 1 5200
box 0 -120 415 525
<< labels >>
rlabel space 4180 7980 4180 7980 7 VPP
rlabel metal3 -120 8705 -120 8705 7 Vref
rlabel space 4195 2500 4195 2500 7 VPP2
rlabel space 170 8545 170 8545 7 Vn
rlabel space 90 8930 90 8930 7 Vp
rlabel locali 15 17275 15 17275 7 Vp
rlabel locali 5025 17935 5025 17935 7 Vref
<< end >>
