magic
tech sky130A
timestamp 1620220727
<< nwell >>
rect -120 350 85 590
<< nmos >>
rect 0 135 15 235
<< pmos >>
rect 0 370 15 570
<< ndiff >>
rect -50 220 0 235
rect -50 150 -35 220
rect -15 150 0 220
rect -50 135 0 150
rect 15 220 65 235
rect 15 150 30 220
rect 50 150 65 220
rect 15 135 65 150
<< pdiff >>
rect -50 555 0 570
rect -50 485 -35 555
rect -15 485 0 555
rect -50 455 0 485
rect -50 385 -35 455
rect -15 385 0 455
rect -50 370 0 385
rect 15 555 65 570
rect 15 485 30 555
rect 50 485 65 555
rect 15 455 65 485
rect 15 385 30 455
rect 50 385 65 455
rect 15 370 65 385
<< ndiffc >>
rect -35 150 -15 220
rect 30 150 50 220
<< pdiffc >>
rect -35 485 -15 555
rect -35 385 -15 455
rect 30 485 50 555
rect 30 385 50 455
<< psubdiff >>
rect -100 220 -50 235
rect -100 150 -85 220
rect -65 150 -50 220
rect -100 135 -50 150
<< nsubdiff >>
rect -100 555 -50 570
rect -100 485 -85 555
rect -65 485 -50 555
rect -100 455 -50 485
rect -100 385 -85 455
rect -65 385 -50 455
rect -100 370 -50 385
<< psubdiffcont >>
rect -85 150 -65 220
<< nsubdiffcont >>
rect -85 485 -65 555
rect -85 385 -65 455
<< poly >>
rect 0 570 15 585
rect 0 235 15 370
rect 0 120 15 135
<< locali >>
rect -95 555 -5 565
rect -95 485 -85 555
rect -65 485 -35 555
rect -15 485 -5 555
rect -95 455 -5 485
rect -95 385 -85 455
rect -65 385 -35 455
rect -15 385 -5 455
rect -95 375 -5 385
rect 20 555 60 565
rect 20 485 30 555
rect 50 485 60 555
rect 20 455 60 485
rect 20 385 30 455
rect 50 385 60 455
rect 20 375 60 385
rect 40 230 60 235
rect -95 220 -5 230
rect -95 150 -85 220
rect -65 150 -35 220
rect -15 150 -5 220
rect -95 140 -5 150
rect 20 220 60 230
rect 20 150 30 220
rect 50 150 60 220
rect 20 140 60 150
<< viali >>
rect -85 485 -65 555
rect -35 485 -15 555
rect -85 385 -65 455
rect -35 385 -15 455
rect -85 150 -65 220
rect -35 150 -15 220
<< metal1 >>
rect -120 555 85 565
rect -120 485 -85 555
rect -65 485 -35 555
rect -15 485 85 555
rect -120 455 85 485
rect -120 385 -85 455
rect -65 385 -35 455
rect -15 385 85 455
rect -120 375 85 385
rect -120 220 85 330
rect -120 150 -85 220
rect -65 150 -35 220
rect -15 150 85 220
rect -120 140 85 150
<< end >>
