magic
tech sky130A
magscale 1 2
timestamp 1620683432
<< nwell >>
rect -410 9300 4130 9800
rect 660 9060 870 9300
rect 2880 9240 3230 9300
rect 2880 9060 3090 9240
rect -410 7750 4130 8150
rect 680 7530 890 7750
rect 2840 7510 3050 7750
rect -410 5880 4130 6280
rect 430 5490 750 5880
rect 2720 5790 3710 5880
rect 2990 5490 3310 5790
<< nmos >>
rect -240 8690 -120 8990
rect 0 8690 120 8990
rect 240 8690 360 8990
rect 480 8690 600 8990
rect 720 8690 840 8990
rect 960 8690 1080 8990
rect 1200 8690 1320 8990
rect 1440 8690 1560 8990
rect 1680 8690 1800 8990
rect 1920 8690 2040 8990
rect 2160 8690 2280 8990
rect 2400 8690 2520 8990
rect 2640 8690 2760 8990
rect 2880 8690 3000 8990
rect 3120 8690 3240 8990
rect 3360 8690 3480 8990
rect 3600 8690 3720 8990
rect 3840 8690 3960 8990
rect -240 6920 -120 7220
rect 0 6920 120 7220
rect 240 6920 360 7220
rect 480 6920 600 7220
rect 720 6920 840 7220
rect 960 6920 1080 7220
rect 1200 6920 1320 7220
rect 1440 6920 1560 7220
rect 1680 6920 1800 7220
rect 1920 6920 2040 7220
rect 2160 6920 2280 7220
rect 2400 6920 2520 7220
rect 2640 6920 2760 7220
rect 2880 6920 3000 7220
rect 3120 6920 3240 7220
rect 3360 6920 3480 7220
rect 3600 6920 3720 7220
rect 3840 6920 3960 7220
rect -240 4860 -120 5160
rect 0 4860 120 5160
rect 240 4860 360 5160
rect 480 4860 600 5160
rect 720 4860 840 5160
rect 960 4860 1080 5160
rect 1200 4860 1320 5160
rect 1440 4860 1560 5160
rect 1680 4860 1800 5160
rect 1920 4860 2040 5160
rect 2160 4860 2280 5160
rect 2400 4860 2520 5160
rect 2640 4860 2760 5160
rect 2880 4860 3000 5160
rect 3120 4860 3240 5160
rect 3360 4860 3480 5160
rect 3600 4860 3720 5160
rect 3840 4860 3960 5160
<< pmos >>
rect -240 9350 -120 9650
rect 0 9350 120 9650
rect 240 9350 360 9650
rect 480 9350 600 9650
rect 720 9350 840 9650
rect 960 9350 1080 9650
rect 1200 9350 1320 9650
rect 1440 9350 1560 9650
rect 1680 9350 1800 9650
rect 1920 9350 2040 9650
rect 2160 9350 2280 9650
rect 2400 9350 2520 9650
rect 2640 9350 2760 9650
rect 2880 9350 3000 9650
rect 3120 9350 3240 9650
rect 3360 9350 3480 9650
rect 3600 9350 3720 9650
rect 3840 9350 3960 9650
rect -240 7800 -120 8100
rect 0 7800 120 8100
rect 240 7800 360 8100
rect 480 7800 600 8100
rect 720 7800 840 8100
rect 960 7800 1080 8100
rect 1200 7800 1320 8100
rect 1440 7800 1560 8100
rect 1680 7800 1800 8100
rect 1920 7800 2040 8100
rect 2160 7800 2280 8100
rect 2400 7800 2520 8100
rect 2640 7800 2760 8100
rect 2880 7800 3000 8100
rect 3120 7800 3240 8100
rect 3360 7800 3480 8100
rect 3600 7800 3720 8100
rect 3840 7800 3960 8100
rect -240 5930 -120 6230
rect 0 5930 120 6230
rect 240 5930 360 6230
rect 480 5930 600 6230
rect 720 5930 840 6230
rect 960 5930 1080 6230
rect 1200 5930 1320 6230
rect 1440 5930 1560 6230
rect 1680 5930 1800 6230
rect 1920 5930 2040 6230
rect 2160 5930 2280 6230
rect 2400 5930 2520 6230
rect 2640 5930 2760 6230
rect 2880 5930 3000 6230
rect 3120 5930 3240 6230
rect 3360 5930 3480 6230
rect 3600 5930 3720 6230
rect 3840 5930 3960 6230
<< ndiff >>
rect -360 8960 -240 8990
rect -360 8720 -330 8960
rect -270 8720 -240 8960
rect -360 8690 -240 8720
rect -120 8960 0 8990
rect -120 8720 -90 8960
rect -30 8720 0 8960
rect -120 8690 0 8720
rect 120 8960 240 8990
rect 120 8720 150 8960
rect 210 8720 240 8960
rect 120 8690 240 8720
rect 360 8960 480 8990
rect 360 8720 390 8960
rect 450 8720 480 8960
rect 360 8690 480 8720
rect 600 8960 720 8990
rect 600 8720 630 8960
rect 690 8720 720 8960
rect 600 8690 720 8720
rect 840 8960 960 8990
rect 840 8720 870 8960
rect 930 8720 960 8960
rect 840 8690 960 8720
rect 1080 8960 1200 8990
rect 1080 8720 1110 8960
rect 1170 8720 1200 8960
rect 1080 8690 1200 8720
rect 1320 8960 1440 8990
rect 1320 8720 1350 8960
rect 1410 8720 1440 8960
rect 1320 8690 1440 8720
rect 1560 8960 1680 8990
rect 1560 8720 1590 8960
rect 1650 8720 1680 8960
rect 1560 8690 1680 8720
rect 1800 8960 1920 8990
rect 1800 8720 1830 8960
rect 1890 8720 1920 8960
rect 1800 8690 1920 8720
rect 2040 8960 2160 8990
rect 2040 8720 2070 8960
rect 2130 8720 2160 8960
rect 2040 8690 2160 8720
rect 2280 8960 2400 8990
rect 2280 8720 2310 8960
rect 2370 8720 2400 8960
rect 2280 8690 2400 8720
rect 2520 8960 2640 8990
rect 2520 8720 2550 8960
rect 2610 8720 2640 8960
rect 2520 8690 2640 8720
rect 2760 8960 2880 8990
rect 2760 8720 2790 8960
rect 2850 8720 2880 8960
rect 2760 8690 2880 8720
rect 3000 8960 3120 8990
rect 3000 8720 3030 8960
rect 3090 8720 3120 8960
rect 3000 8690 3120 8720
rect 3240 8960 3360 8990
rect 3240 8720 3270 8960
rect 3330 8720 3360 8960
rect 3240 8690 3360 8720
rect 3480 8960 3600 8990
rect 3480 8720 3510 8960
rect 3570 8720 3600 8960
rect 3480 8690 3600 8720
rect 3720 8960 3840 8990
rect 3720 8720 3750 8960
rect 3810 8720 3840 8960
rect 3720 8690 3840 8720
rect 3960 8960 4080 8990
rect 3960 8720 3990 8960
rect 4050 8720 4080 8960
rect 3960 8690 4080 8720
rect -360 7190 -240 7220
rect -360 6950 -330 7190
rect -270 6950 -240 7190
rect -360 6920 -240 6950
rect -120 7190 0 7220
rect -120 6950 -90 7190
rect -30 6950 0 7190
rect -120 6920 0 6950
rect 120 7190 240 7220
rect 120 6950 150 7190
rect 210 6950 240 7190
rect 120 6920 240 6950
rect 360 7190 480 7220
rect 360 6950 390 7190
rect 450 6950 480 7190
rect 360 6920 480 6950
rect 600 7190 720 7220
rect 600 6950 630 7190
rect 690 6950 720 7190
rect 600 6920 720 6950
rect 840 7190 960 7220
rect 840 6950 870 7190
rect 930 6950 960 7190
rect 840 6920 960 6950
rect 1080 7190 1200 7220
rect 1080 6950 1110 7190
rect 1170 6950 1200 7190
rect 1080 6920 1200 6950
rect 1320 7190 1440 7220
rect 1320 6950 1350 7190
rect 1410 6950 1440 7190
rect 1320 6920 1440 6950
rect 1560 7190 1680 7220
rect 1560 6950 1590 7190
rect 1650 6950 1680 7190
rect 1560 6920 1680 6950
rect 1800 7190 1920 7220
rect 1800 6950 1830 7190
rect 1890 6950 1920 7190
rect 1800 6920 1920 6950
rect 2040 7190 2160 7220
rect 2040 6950 2070 7190
rect 2130 6950 2160 7190
rect 2040 6920 2160 6950
rect 2280 7190 2400 7220
rect 2280 6950 2310 7190
rect 2370 6950 2400 7190
rect 2280 6920 2400 6950
rect 2520 7190 2640 7220
rect 2520 6950 2550 7190
rect 2610 6950 2640 7190
rect 2520 6920 2640 6950
rect 2760 7190 2880 7220
rect 2760 6950 2790 7190
rect 2850 6950 2880 7190
rect 2760 6920 2880 6950
rect 3000 7190 3120 7220
rect 3000 6950 3030 7190
rect 3090 6950 3120 7190
rect 3000 6920 3120 6950
rect 3240 7190 3360 7220
rect 3240 6950 3270 7190
rect 3330 6950 3360 7190
rect 3240 6920 3360 6950
rect 3480 7190 3600 7220
rect 3480 6950 3510 7190
rect 3570 6950 3600 7190
rect 3480 6920 3600 6950
rect 3720 7190 3840 7220
rect 3720 6950 3750 7190
rect 3810 6950 3840 7190
rect 3720 6920 3840 6950
rect 3960 7190 4080 7220
rect 3960 6950 3990 7190
rect 4050 6950 4080 7190
rect 3960 6920 4080 6950
rect -360 5130 -240 5160
rect -360 4890 -330 5130
rect -270 4890 -240 5130
rect -360 4860 -240 4890
rect -120 5130 0 5160
rect -120 4890 -90 5130
rect -30 4890 0 5130
rect -120 4860 0 4890
rect 120 5130 240 5160
rect 120 4890 150 5130
rect 210 4890 240 5130
rect 120 4860 240 4890
rect 360 5130 480 5160
rect 360 4890 390 5130
rect 450 4890 480 5130
rect 360 4860 480 4890
rect 600 5130 720 5160
rect 600 4890 630 5130
rect 690 4890 720 5130
rect 600 4860 720 4890
rect 840 5130 960 5160
rect 840 4890 870 5130
rect 930 4890 960 5130
rect 840 4860 960 4890
rect 1080 5130 1200 5160
rect 1080 4890 1110 5130
rect 1170 4890 1200 5130
rect 1080 4860 1200 4890
rect 1320 5130 1440 5160
rect 1320 4890 1350 5130
rect 1410 4890 1440 5130
rect 1320 4860 1440 4890
rect 1560 5130 1680 5160
rect 1560 4890 1590 5130
rect 1650 4890 1680 5130
rect 1560 4860 1680 4890
rect 1800 5130 1920 5160
rect 1800 4890 1830 5130
rect 1890 4890 1920 5130
rect 1800 4860 1920 4890
rect 2040 5130 2160 5160
rect 2040 4890 2070 5130
rect 2130 4890 2160 5130
rect 2040 4860 2160 4890
rect 2280 5130 2400 5160
rect 2280 4890 2310 5130
rect 2370 4890 2400 5130
rect 2280 4860 2400 4890
rect 2520 5130 2640 5160
rect 2520 4890 2550 5130
rect 2610 4890 2640 5130
rect 2520 4860 2640 4890
rect 2760 5130 2880 5160
rect 2760 4890 2790 5130
rect 2850 4890 2880 5130
rect 2760 4860 2880 4890
rect 3000 5130 3120 5160
rect 3000 4890 3030 5130
rect 3090 4890 3120 5130
rect 3000 4860 3120 4890
rect 3240 5130 3360 5160
rect 3240 4890 3270 5130
rect 3330 4890 3360 5130
rect 3240 4860 3360 4890
rect 3480 5130 3600 5160
rect 3480 4890 3510 5130
rect 3570 4890 3600 5130
rect 3480 4860 3600 4890
rect 3720 5130 3840 5160
rect 3720 4890 3750 5130
rect 3810 4890 3840 5130
rect 3720 4860 3840 4890
rect 3960 5130 4080 5160
rect 3960 4890 3990 5130
rect 4050 4890 4080 5130
rect 3960 4860 4080 4890
<< pdiff >>
rect -360 9620 -240 9650
rect -360 9380 -330 9620
rect -270 9380 -240 9620
rect -360 9350 -240 9380
rect -120 9620 0 9650
rect -120 9380 -90 9620
rect -30 9380 0 9620
rect -120 9350 0 9380
rect 120 9620 240 9650
rect 120 9380 150 9620
rect 210 9380 240 9620
rect 120 9350 240 9380
rect 360 9620 480 9650
rect 360 9380 390 9620
rect 450 9380 480 9620
rect 360 9350 480 9380
rect 600 9620 720 9650
rect 600 9380 630 9620
rect 690 9380 720 9620
rect 600 9350 720 9380
rect 840 9620 960 9650
rect 840 9380 870 9620
rect 930 9380 960 9620
rect 840 9350 960 9380
rect 1080 9620 1200 9650
rect 1080 9380 1110 9620
rect 1170 9380 1200 9620
rect 1080 9350 1200 9380
rect 1320 9620 1440 9650
rect 1320 9380 1350 9620
rect 1410 9380 1440 9620
rect 1320 9350 1440 9380
rect 1560 9620 1680 9650
rect 1560 9380 1590 9620
rect 1650 9380 1680 9620
rect 1560 9350 1680 9380
rect 1800 9620 1920 9650
rect 1800 9380 1830 9620
rect 1890 9380 1920 9620
rect 1800 9350 1920 9380
rect 2040 9620 2160 9650
rect 2040 9380 2070 9620
rect 2130 9380 2160 9620
rect 2040 9350 2160 9380
rect 2280 9620 2400 9650
rect 2280 9380 2310 9620
rect 2370 9380 2400 9620
rect 2280 9350 2400 9380
rect 2520 9620 2640 9650
rect 2520 9380 2550 9620
rect 2610 9380 2640 9620
rect 2520 9350 2640 9380
rect 2760 9620 2880 9650
rect 2760 9380 2790 9620
rect 2850 9380 2880 9620
rect 2760 9350 2880 9380
rect 3000 9620 3120 9650
rect 3000 9380 3030 9620
rect 3090 9380 3120 9620
rect 3000 9350 3120 9380
rect 3240 9620 3360 9650
rect 3240 9380 3270 9620
rect 3330 9380 3360 9620
rect 3240 9350 3360 9380
rect 3480 9620 3600 9650
rect 3480 9380 3510 9620
rect 3570 9380 3600 9620
rect 3480 9350 3600 9380
rect 3720 9620 3840 9650
rect 3720 9380 3750 9620
rect 3810 9380 3840 9620
rect 3720 9350 3840 9380
rect 3960 9620 4080 9650
rect 3960 9380 3990 9620
rect 4050 9380 4080 9620
rect 3960 9350 4080 9380
rect -360 8070 -240 8100
rect -360 7830 -330 8070
rect -270 7830 -240 8070
rect -360 7800 -240 7830
rect -120 8070 0 8100
rect -120 7830 -90 8070
rect -30 7830 0 8070
rect -120 7800 0 7830
rect 120 8070 240 8100
rect 120 7830 150 8070
rect 210 7830 240 8070
rect 120 7800 240 7830
rect 360 8070 480 8100
rect 360 7830 390 8070
rect 450 7830 480 8070
rect 360 7800 480 7830
rect 600 8070 720 8100
rect 600 7830 630 8070
rect 690 7830 720 8070
rect 600 7800 720 7830
rect 840 8070 960 8100
rect 840 7830 870 8070
rect 930 7830 960 8070
rect 840 7800 960 7830
rect 1080 8070 1200 8100
rect 1080 7830 1110 8070
rect 1170 7830 1200 8070
rect 1080 7800 1200 7830
rect 1320 8070 1440 8100
rect 1320 7830 1350 8070
rect 1410 7830 1440 8070
rect 1320 7800 1440 7830
rect 1560 8070 1680 8100
rect 1560 7830 1590 8070
rect 1650 7830 1680 8070
rect 1560 7800 1680 7830
rect 1800 8070 1920 8100
rect 1800 7830 1830 8070
rect 1890 7830 1920 8070
rect 1800 7800 1920 7830
rect 2040 8070 2160 8100
rect 2040 7830 2070 8070
rect 2130 7830 2160 8070
rect 2040 7800 2160 7830
rect 2280 8070 2400 8100
rect 2280 7830 2310 8070
rect 2370 7830 2400 8070
rect 2280 7800 2400 7830
rect 2520 8070 2640 8100
rect 2520 7830 2550 8070
rect 2610 7830 2640 8070
rect 2520 7800 2640 7830
rect 2760 8070 2880 8100
rect 2760 7830 2790 8070
rect 2850 7830 2880 8070
rect 2760 7800 2880 7830
rect 3000 8070 3120 8100
rect 3000 7830 3030 8070
rect 3090 7830 3120 8070
rect 3000 7800 3120 7830
rect 3240 8070 3360 8100
rect 3240 7830 3270 8070
rect 3330 7830 3360 8070
rect 3240 7800 3360 7830
rect 3480 8070 3600 8100
rect 3480 7830 3510 8070
rect 3570 7830 3600 8070
rect 3480 7800 3600 7830
rect 3720 8070 3840 8100
rect 3720 7830 3750 8070
rect 3810 7830 3840 8070
rect 3720 7800 3840 7830
rect 3960 8070 4080 8100
rect 3960 7830 3990 8070
rect 4050 7830 4080 8070
rect 3960 7800 4080 7830
rect -360 6200 -240 6230
rect -360 5960 -330 6200
rect -270 5960 -240 6200
rect -360 5930 -240 5960
rect -120 6200 0 6230
rect -120 5960 -90 6200
rect -30 5960 0 6200
rect -120 5930 0 5960
rect 120 6200 240 6230
rect 120 5960 150 6200
rect 210 5960 240 6200
rect 120 5930 240 5960
rect 360 6200 480 6230
rect 360 5960 390 6200
rect 450 5960 480 6200
rect 360 5930 480 5960
rect 600 6200 720 6230
rect 600 5960 630 6200
rect 690 5960 720 6200
rect 600 5930 720 5960
rect 840 6200 960 6230
rect 840 5960 870 6200
rect 930 5960 960 6200
rect 840 5930 960 5960
rect 1080 6200 1200 6230
rect 1080 5960 1110 6200
rect 1170 5960 1200 6200
rect 1080 5930 1200 5960
rect 1320 6200 1440 6230
rect 1320 5960 1350 6200
rect 1410 5960 1440 6200
rect 1320 5930 1440 5960
rect 1560 6200 1680 6230
rect 1560 5960 1590 6200
rect 1650 5960 1680 6200
rect 1560 5930 1680 5960
rect 1800 6200 1920 6230
rect 1800 5960 1830 6200
rect 1890 5960 1920 6200
rect 1800 5930 1920 5960
rect 2040 6200 2160 6230
rect 2040 5960 2070 6200
rect 2130 5960 2160 6200
rect 2040 5930 2160 5960
rect 2280 6200 2400 6230
rect 2280 5960 2310 6200
rect 2370 5960 2400 6200
rect 2280 5930 2400 5960
rect 2520 6200 2640 6230
rect 2520 5960 2550 6200
rect 2610 5960 2640 6200
rect 2520 5930 2640 5960
rect 2760 6200 2880 6230
rect 2760 5960 2790 6200
rect 2850 5960 2880 6200
rect 2760 5930 2880 5960
rect 3000 6200 3120 6230
rect 3000 5960 3030 6200
rect 3090 5960 3120 6200
rect 3000 5930 3120 5960
rect 3240 6200 3360 6230
rect 3240 5960 3270 6200
rect 3330 5960 3360 6200
rect 3240 5930 3360 5960
rect 3480 6200 3600 6230
rect 3480 5960 3510 6200
rect 3570 5960 3600 6200
rect 3480 5930 3600 5960
rect 3720 6200 3840 6230
rect 3720 5960 3750 6200
rect 3810 5960 3840 6200
rect 3720 5930 3840 5960
rect 3960 6200 4080 6230
rect 3960 5960 3990 6200
rect 4050 5960 4080 6200
rect 3960 5930 4080 5960
<< ndiffc >>
rect -330 8720 -270 8960
rect -90 8720 -30 8960
rect 150 8720 210 8960
rect 390 8720 450 8960
rect 630 8720 690 8960
rect 870 8720 930 8960
rect 1110 8720 1170 8960
rect 1350 8720 1410 8960
rect 1590 8720 1650 8960
rect 1830 8720 1890 8960
rect 2070 8720 2130 8960
rect 2310 8720 2370 8960
rect 2550 8720 2610 8960
rect 2790 8720 2850 8960
rect 3030 8720 3090 8960
rect 3270 8720 3330 8960
rect 3510 8720 3570 8960
rect 3750 8720 3810 8960
rect 3990 8720 4050 8960
rect -330 6950 -270 7190
rect -90 6950 -30 7190
rect 150 6950 210 7190
rect 390 6950 450 7190
rect 630 6950 690 7190
rect 870 6950 930 7190
rect 1110 6950 1170 7190
rect 1350 6950 1410 7190
rect 1590 6950 1650 7190
rect 1830 6950 1890 7190
rect 2070 6950 2130 7190
rect 2310 6950 2370 7190
rect 2550 6950 2610 7190
rect 2790 6950 2850 7190
rect 3030 6950 3090 7190
rect 3270 6950 3330 7190
rect 3510 6950 3570 7190
rect 3750 6950 3810 7190
rect 3990 6950 4050 7190
rect -330 4890 -270 5130
rect -90 4890 -30 5130
rect 150 4890 210 5130
rect 390 4890 450 5130
rect 630 4890 690 5130
rect 870 4890 930 5130
rect 1110 4890 1170 5130
rect 1350 4890 1410 5130
rect 1590 4890 1650 5130
rect 1830 4890 1890 5130
rect 2070 4890 2130 5130
rect 2310 4890 2370 5130
rect 2550 4890 2610 5130
rect 2790 4890 2850 5130
rect 3030 4890 3090 5130
rect 3270 4890 3330 5130
rect 3510 4890 3570 5130
rect 3750 4890 3810 5130
rect 3990 4890 4050 5130
<< pdiffc >>
rect -330 9380 -270 9620
rect -90 9380 -30 9620
rect 150 9380 210 9620
rect 390 9380 450 9620
rect 630 9380 690 9620
rect 870 9380 930 9620
rect 1110 9380 1170 9620
rect 1350 9380 1410 9620
rect 1590 9380 1650 9620
rect 1830 9380 1890 9620
rect 2070 9380 2130 9620
rect 2310 9380 2370 9620
rect 2550 9380 2610 9620
rect 2790 9380 2850 9620
rect 3030 9380 3090 9620
rect 3270 9380 3330 9620
rect 3510 9380 3570 9620
rect 3750 9380 3810 9620
rect 3990 9380 4050 9620
rect -330 7830 -270 8070
rect -90 7830 -30 8070
rect 150 7830 210 8070
rect 390 7830 450 8070
rect 630 7830 690 8070
rect 870 7830 930 8070
rect 1110 7830 1170 8070
rect 1350 7830 1410 8070
rect 1590 7830 1650 8070
rect 1830 7830 1890 8070
rect 2070 7830 2130 8070
rect 2310 7830 2370 8070
rect 2550 7830 2610 8070
rect 2790 7830 2850 8070
rect 3030 7830 3090 8070
rect 3270 7830 3330 8070
rect 3510 7830 3570 8070
rect 3750 7830 3810 8070
rect 3990 7830 4050 8070
rect -330 5960 -270 6200
rect -90 5960 -30 6200
rect 150 5960 210 6200
rect 390 5960 450 6200
rect 630 5960 690 6200
rect 870 5960 930 6200
rect 1110 5960 1170 6200
rect 1350 5960 1410 6200
rect 1590 5960 1650 6200
rect 1830 5960 1890 6200
rect 2070 5960 2130 6200
rect 2310 5960 2370 6200
rect 2550 5960 2610 6200
rect 2790 5960 2850 6200
rect 3030 5960 3090 6200
rect 3270 5960 3330 6200
rect 3510 5960 3570 6200
rect 3750 5960 3810 6200
rect 3990 5960 4050 6200
<< psubdiff >>
rect 330 9150 450 9180
rect 330 9090 360 9150
rect 420 9090 450 9150
rect 330 9060 450 9090
rect 3440 9180 3560 9210
rect 3440 9120 3470 9180
rect 3530 9120 3560 9180
rect 3440 9090 3560 9120
rect 330 7510 450 7540
rect 330 7440 360 7510
rect 420 7440 450 7510
rect 330 7410 450 7440
rect 3350 7490 3470 7520
rect 3350 7420 3380 7490
rect 3440 7420 3470 7490
rect 3350 7390 3470 7420
rect 900 5460 1140 5490
rect 900 5280 930 5460
rect 1110 5280 1140 5460
rect 2580 5460 2820 5490
rect 900 5250 1140 5280
rect 2580 5280 2610 5460
rect 2790 5280 2820 5460
rect 2580 5250 2820 5280
<< nsubdiff >>
rect 700 9190 820 9210
rect 700 9130 730 9190
rect 790 9130 820 9190
rect 700 9100 820 9130
rect 2920 9190 3040 9210
rect 2920 9130 2950 9190
rect 3010 9130 3040 9190
rect 2920 9100 3040 9130
rect 720 7670 840 7700
rect 720 7600 750 7670
rect 810 7600 840 7670
rect 2880 7650 3000 7680
rect 720 7570 840 7600
rect 2880 7580 2910 7650
rect 2970 7580 3000 7650
rect 2880 7550 3000 7580
rect 470 5740 710 5770
rect 470 5560 500 5740
rect 680 5560 710 5740
rect 3030 5740 3270 5770
rect 470 5530 710 5560
rect 3030 5560 3060 5740
rect 3240 5560 3270 5740
rect 3030 5530 3270 5560
<< psubdiffcont >>
rect 360 9090 420 9150
rect 3470 9120 3530 9180
rect 360 7440 420 7510
rect 3380 7420 3440 7490
rect 930 5280 1110 5460
rect 2610 5280 2790 5460
<< nsubdiffcont >>
rect 730 9130 790 9190
rect 2950 9130 3010 9190
rect 750 7600 810 7670
rect 2910 7580 2970 7650
rect 500 5560 680 5740
rect 3060 5560 3240 5740
<< poly >>
rect -500 9830 2760 9860
rect -240 9650 -120 9680
rect 0 9650 120 9680
rect 240 9650 360 9680
rect 480 9650 600 9680
rect 720 9650 840 9680
rect 960 9650 1080 9830
rect 1200 9750 1320 9780
rect 1200 9710 1250 9750
rect 1290 9710 1320 9750
rect 1200 9650 1320 9710
rect 1440 9730 2280 9770
rect 1440 9650 1560 9730
rect 1680 9650 1800 9680
rect 1920 9650 2040 9680
rect 2160 9650 2280 9730
rect 2400 9750 2520 9780
rect 2400 9710 2430 9750
rect 2470 9710 2520 9750
rect 2400 9650 2520 9710
rect 2640 9650 2760 9830
rect 2880 9650 3000 9680
rect 3120 9650 3240 9680
rect 3360 9650 3480 9680
rect 3600 9650 3720 9680
rect 3840 9650 3960 9680
rect -240 9320 -120 9350
rect 0 9320 120 9350
rect 240 9320 360 9350
rect 480 9320 600 9350
rect 720 9320 840 9350
rect -350 9300 840 9320
rect -350 9260 -330 9300
rect -140 9260 -90 9300
rect 100 9260 150 9300
rect 340 9260 390 9300
rect 580 9260 630 9300
rect 820 9260 840 9300
rect -350 9240 840 9260
rect -240 8990 -120 9020
rect 0 8990 120 9020
rect 240 8990 360 9020
rect 480 8990 600 9020
rect 720 8990 840 9020
rect 960 8990 1080 9350
rect 1200 9320 1320 9350
rect 1440 9270 1560 9350
rect 1200 9240 1560 9270
rect 1200 8990 1320 9240
rect 1680 9180 1800 9350
rect 1920 9180 2040 9350
rect 2160 9270 2280 9350
rect 2400 9320 2520 9350
rect 2160 9240 2520 9270
rect 1680 9160 2040 9180
rect 1680 9150 1840 9160
rect 1820 9120 1840 9150
rect 1880 9150 2040 9160
rect 1880 9120 1900 9150
rect 1820 9100 1900 9120
rect 1440 8990 1560 9020
rect 1680 8990 1800 9020
rect 1920 8990 2040 9020
rect 2160 8990 2280 9020
rect 2400 8990 2520 9240
rect 2640 8990 2760 9350
rect 2880 9320 3000 9350
rect 3120 9320 3240 9350
rect 3360 9320 3480 9350
rect 3600 9320 3720 9350
rect 3840 9320 3960 9350
rect 2880 9300 4070 9320
rect 2880 9260 2900 9300
rect 3090 9260 3140 9300
rect 3330 9260 3380 9300
rect 3570 9260 3620 9300
rect 3810 9260 3860 9300
rect 4050 9260 4070 9300
rect 2880 9240 4070 9260
rect 4040 9080 4120 9100
rect 4040 9040 4060 9080
rect 4100 9050 4120 9080
rect 4100 9040 4150 9050
rect 4040 9020 4150 9040
rect 2880 8990 3000 9020
rect 3120 8990 3240 9020
rect 3360 8990 3480 9020
rect 3600 8990 3720 9020
rect 3840 8990 3960 9020
rect -240 8660 -120 8690
rect 0 8660 120 8690
rect 240 8660 360 8690
rect 480 8660 600 8690
rect 720 8660 840 8690
rect 960 8660 1080 8690
rect -350 8640 840 8660
rect -350 8600 -330 8640
rect -140 8600 -90 8640
rect 100 8600 150 8640
rect 340 8600 390 8640
rect 580 8600 630 8640
rect 820 8600 840 8640
rect -350 8580 840 8600
rect 1200 8410 1320 8690
rect 1440 8660 1560 8690
rect 1450 8650 1530 8660
rect 1450 8610 1470 8650
rect 1510 8610 1530 8650
rect 1450 8590 1530 8610
rect 1680 8610 1800 8690
rect 1920 8610 2040 8690
rect 2160 8660 2280 8690
rect 2400 8660 2520 8690
rect 2640 8660 2760 8690
rect 2880 8660 3000 8690
rect 3120 8660 3240 8690
rect 3360 8660 3480 8690
rect 3600 8660 3720 8690
rect 3840 8660 3960 8690
rect -500 8380 1320 8410
rect 1680 8580 2040 8610
rect 2190 8650 2270 8660
rect 2190 8610 2210 8650
rect 2250 8610 2270 8650
rect 2190 8590 2270 8610
rect 2880 8640 4070 8660
rect 2880 8600 2900 8640
rect 3090 8600 3140 8640
rect 3330 8600 3380 8640
rect 3570 8600 3620 8640
rect 3810 8600 3860 8640
rect 4050 8600 4070 8640
rect 2880 8580 4070 8600
rect 1680 8330 1710 8580
rect -440 8300 1710 8330
rect -440 7380 -410 8300
rect 4120 8210 4150 9020
rect 720 8180 4150 8210
rect -240 8100 -120 8130
rect 0 8100 120 8130
rect 240 8100 360 8130
rect 480 8100 600 8130
rect 720 8100 840 8180
rect 960 8100 1080 8130
rect 1200 8100 1320 8130
rect 1440 8100 1560 8180
rect 1680 8100 1800 8130
rect 1920 8100 2040 8130
rect 2160 8100 2280 8180
rect 2400 8100 2520 8130
rect 2640 8100 2760 8130
rect 2880 8100 3000 8180
rect 3120 8100 3240 8130
rect 3360 8100 3480 8130
rect 3600 8100 3720 8130
rect 3840 8100 3960 8130
rect -240 7770 -120 7800
rect 0 7770 120 7800
rect 240 7770 360 7800
rect 480 7770 600 7800
rect 720 7770 840 7800
rect -350 7750 600 7770
rect -350 7710 -330 7750
rect -140 7710 -90 7750
rect 100 7710 150 7750
rect 340 7710 390 7750
rect 580 7710 600 7750
rect -350 7690 600 7710
rect 960 7750 1080 7800
rect 1200 7770 1320 7800
rect 1440 7770 1560 7800
rect 960 7710 980 7750
rect 1060 7710 1080 7750
rect 960 7690 1080 7710
rect 1240 7750 1320 7770
rect 1240 7710 1260 7750
rect 1300 7710 1320 7750
rect 1240 7690 1320 7710
rect 1680 7750 1800 7800
rect 1680 7710 1700 7750
rect 1780 7710 1800 7750
rect 1680 7690 1800 7710
rect 1920 7750 2040 7800
rect 2160 7770 2280 7800
rect 2400 7770 2520 7800
rect 1920 7710 1940 7750
rect 2020 7710 2040 7750
rect 1920 7690 2040 7710
rect 2400 7750 2480 7770
rect 2400 7710 2420 7750
rect 2460 7710 2480 7750
rect 2400 7690 2480 7710
rect 2640 7750 2760 7800
rect 2880 7770 3000 7800
rect 3120 7770 3240 7800
rect 3360 7770 3480 7800
rect 3600 7770 3720 7800
rect 3840 7770 3960 7800
rect 2640 7710 2660 7750
rect 2740 7710 2760 7750
rect 2640 7690 2760 7710
rect 3120 7750 4070 7770
rect 3120 7710 3140 7750
rect 3330 7710 3380 7750
rect 3570 7710 3620 7750
rect 3810 7710 3860 7750
rect 4050 7710 4070 7750
rect 3120 7690 4070 7710
rect 1820 7630 1900 7650
rect 1820 7590 1840 7630
rect 1880 7590 1900 7630
rect 1820 7570 1900 7590
rect 1840 7450 1880 7570
rect 3200 7550 3560 7590
rect 3200 7450 3240 7550
rect 1820 7430 3240 7450
rect 1820 7390 1840 7430
rect 1880 7410 3240 7430
rect 3520 7510 3560 7550
rect 3520 7490 4070 7510
rect 3520 7470 4010 7490
rect 3990 7450 4010 7470
rect 4050 7450 4070 7490
rect 3990 7430 4070 7450
rect 1880 7390 1900 7410
rect -440 7350 840 7380
rect 1820 7370 1900 7390
rect -240 7220 -120 7250
rect 0 7220 120 7250
rect 240 7220 360 7250
rect 480 7220 600 7250
rect 720 7220 840 7350
rect 960 7310 1080 7330
rect 960 7270 980 7310
rect 1060 7270 1080 7310
rect 960 7220 1080 7270
rect 1240 7310 1320 7330
rect 1240 7270 1260 7310
rect 1300 7270 1320 7310
rect 1240 7250 1320 7270
rect 1680 7310 1800 7330
rect 1680 7270 1700 7310
rect 1780 7270 1800 7310
rect 1200 7220 1320 7250
rect 1440 7220 1560 7250
rect 1680 7220 1800 7270
rect 1920 7310 2040 7330
rect 1920 7270 1940 7310
rect 2020 7270 2040 7310
rect 1920 7220 2040 7270
rect 2400 7310 2480 7330
rect 2400 7270 2420 7310
rect 2460 7270 2480 7310
rect 2400 7250 2480 7270
rect 2640 7310 2760 7330
rect 2640 7270 2660 7310
rect 2740 7270 2760 7310
rect 2160 7220 2280 7250
rect 2400 7220 2520 7250
rect 2640 7220 2760 7270
rect 2880 7220 3000 7250
rect 3120 7220 3240 7250
rect 3360 7220 3480 7250
rect 3600 7220 3720 7250
rect 3840 7220 3960 7250
rect -240 6890 -120 6920
rect 0 6890 120 6920
rect 240 6890 360 6920
rect 480 6890 600 6920
rect -350 6870 600 6890
rect -350 6830 -330 6870
rect -140 6830 -90 6870
rect 100 6830 150 6870
rect 340 6830 390 6870
rect 580 6830 600 6870
rect -350 6810 600 6830
rect 720 6840 840 6920
rect 960 6890 1080 6920
rect 1200 6890 1320 6920
rect 1440 6840 1560 6920
rect 1680 6890 1800 6920
rect 1920 6890 2040 6920
rect 2160 6840 2280 6920
rect 2400 6890 2520 6920
rect 2640 6890 2760 6920
rect 2880 6840 3000 6920
rect 720 6810 3000 6840
rect 3120 6890 3240 6920
rect 3360 6890 3480 6920
rect 3600 6890 3720 6920
rect 3840 6890 3960 6920
rect 3120 6870 4070 6890
rect 3120 6830 3140 6870
rect 3330 6830 3380 6870
rect 3570 6830 3620 6870
rect 3810 6830 3860 6870
rect 4050 6830 4070 6870
rect 3120 6810 4070 6830
rect 880 6380 920 6810
rect 720 6360 800 6380
rect 720 6320 740 6360
rect 780 6320 800 6360
rect 720 6260 800 6320
rect 860 6360 940 6380
rect 860 6320 880 6360
rect 920 6320 940 6360
rect 860 6300 940 6320
rect 1440 6360 1520 6380
rect 1440 6320 1460 6360
rect 1500 6320 1520 6360
rect 1440 6260 1520 6320
rect 2200 6360 2280 6380
rect 2200 6320 2220 6360
rect 2260 6320 2280 6360
rect 2200 6260 2280 6320
rect 2920 6360 3000 6380
rect 2920 6320 2940 6360
rect 2980 6320 3000 6360
rect 4120 6350 4150 8180
rect 4300 6440 4380 6460
rect 4300 6400 4320 6440
rect 4360 6400 4380 6440
rect 4300 6380 4380 6400
rect 2920 6260 3000 6320
rect 3600 6320 4150 6350
rect -240 6230 -120 6260
rect 0 6230 120 6260
rect 240 6230 360 6260
rect 480 6230 600 6260
rect 720 6230 840 6260
rect 960 6230 1080 6260
rect 1200 6230 1320 6260
rect 1440 6230 1560 6260
rect 1680 6230 1800 6260
rect 1920 6230 2040 6260
rect 2160 6230 2280 6260
rect 2400 6230 2520 6260
rect 2640 6230 2760 6260
rect 2880 6230 3000 6260
rect 3120 6230 3240 6260
rect 3360 6230 3480 6260
rect 3600 6230 3720 6320
rect 4350 6300 4380 6380
rect 3840 6230 3960 6260
rect -240 5900 -120 5930
rect -350 5880 -120 5900
rect -350 5840 -330 5880
rect -140 5840 -120 5880
rect -350 5820 -120 5840
rect 0 5850 120 5930
rect 240 5850 360 5930
rect 480 5850 600 5930
rect 720 5900 840 5930
rect 960 5850 1080 5930
rect 1200 5850 1320 5930
rect 1440 5900 1560 5930
rect 1680 5850 1800 5930
rect 1920 5850 2040 5930
rect 2160 5900 2280 5930
rect 2400 5850 2520 5930
rect 2640 5850 2760 5930
rect 2880 5900 3000 5930
rect 3120 5850 3240 5930
rect 3360 5850 3480 5930
rect 3600 5850 3720 5930
rect 0 5830 3720 5850
rect 0 5820 1840 5830
rect 1820 5790 1840 5820
rect 1880 5820 3720 5830
rect 3840 5900 3960 5930
rect 3840 5880 4070 5900
rect 3840 5840 3860 5880
rect 4050 5840 4070 5880
rect 3840 5820 4070 5840
rect 1880 5790 1900 5820
rect 1820 5770 1900 5790
rect 1570 5750 1670 5770
rect 1570 5700 1590 5750
rect 1650 5710 1670 5750
rect 2050 5750 2150 5770
rect 2050 5710 2070 5750
rect 1650 5700 2070 5710
rect 2130 5700 2150 5750
rect 850 5670 950 5700
rect 1570 5680 2150 5700
rect 850 5620 870 5670
rect 930 5630 950 5670
rect 2770 5670 2870 5700
rect 2770 5630 2790 5670
rect 930 5620 2790 5630
rect 2850 5620 2870 5670
rect 850 5600 2870 5620
rect 1840 5330 1880 5600
rect 1810 5310 1910 5330
rect 720 5240 840 5280
rect 720 5200 760 5240
rect 800 5200 840 5240
rect -240 5160 -120 5190
rect 0 5160 120 5190
rect 240 5160 360 5190
rect 480 5160 600 5190
rect 720 5160 840 5200
rect 1440 5240 1560 5280
rect 1810 5260 1830 5310
rect 1890 5260 1910 5310
rect 1810 5240 1910 5260
rect 2160 5240 2280 5280
rect 2880 5270 3000 5310
rect 1440 5200 1480 5240
rect 1520 5200 1560 5240
rect 960 5160 1080 5190
rect 1200 5160 1320 5190
rect 1440 5160 1560 5200
rect 2160 5200 2200 5240
rect 2240 5200 2280 5240
rect 1680 5160 1800 5190
rect 1920 5160 2040 5190
rect 2160 5160 2280 5200
rect 2880 5230 2920 5270
rect 2960 5230 3000 5270
rect 2400 5160 2520 5190
rect 2640 5160 2760 5190
rect 2880 5160 3000 5230
rect 3120 5160 3240 5190
rect 3360 5160 3480 5190
rect 3600 5160 3720 5190
rect 3840 5160 3960 5190
rect -240 4830 -120 4860
rect -350 4810 -120 4830
rect -350 4770 -330 4810
rect -140 4770 -120 4810
rect -350 4750 -120 4770
rect 0 4780 120 4860
rect 240 4780 360 4860
rect 480 4780 600 4860
rect 720 4830 840 4860
rect 960 4780 1080 4860
rect 1200 4780 1320 4860
rect 1440 4830 1560 4860
rect 1680 4790 1800 4860
rect 1920 4790 2040 4860
rect 2160 4830 2280 4860
rect 1680 4780 2040 4790
rect 2400 4780 2520 4860
rect 2640 4780 2760 4860
rect 2880 4830 3000 4860
rect 3120 4780 3240 4860
rect 3360 4780 3480 4860
rect 3600 4780 3720 4860
rect 0 4770 3720 4780
rect 0 4750 1840 4770
rect 1820 4730 1840 4750
rect 1880 4750 3720 4770
rect 3840 4830 3960 4860
rect 3840 4810 4070 4830
rect 3840 4770 3860 4810
rect 4050 4770 4070 4810
rect 3840 4750 4070 4770
rect 1880 4730 1900 4750
rect 1820 4710 1900 4730
<< polycont >>
rect 1250 9710 1290 9750
rect 2430 9710 2470 9750
rect -330 9260 -140 9300
rect -90 9260 100 9300
rect 150 9260 340 9300
rect 390 9260 580 9300
rect 630 9260 820 9300
rect 1840 9120 1880 9160
rect 2900 9260 3090 9300
rect 3140 9260 3330 9300
rect 3380 9260 3570 9300
rect 3620 9260 3810 9300
rect 3860 9260 4050 9300
rect 4060 9040 4100 9080
rect -330 8600 -140 8640
rect -90 8600 100 8640
rect 150 8600 340 8640
rect 390 8600 580 8640
rect 630 8600 820 8640
rect 1470 8610 1510 8650
rect 2210 8610 2250 8650
rect 2900 8600 3090 8640
rect 3140 8600 3330 8640
rect 3380 8600 3570 8640
rect 3620 8600 3810 8640
rect 3860 8600 4050 8640
rect -330 7710 -140 7750
rect -90 7710 100 7750
rect 150 7710 340 7750
rect 390 7710 580 7750
rect 980 7710 1060 7750
rect 1260 7710 1300 7750
rect 1700 7710 1780 7750
rect 1940 7710 2020 7750
rect 2420 7710 2460 7750
rect 2660 7710 2740 7750
rect 3140 7710 3330 7750
rect 3380 7710 3570 7750
rect 3620 7710 3810 7750
rect 3860 7710 4050 7750
rect 1840 7590 1880 7630
rect 1840 7390 1880 7430
rect 4010 7450 4050 7490
rect 980 7270 1060 7310
rect 1260 7270 1300 7310
rect 1700 7270 1780 7310
rect 1940 7270 2020 7310
rect 2420 7270 2460 7310
rect 2660 7270 2740 7310
rect -330 6830 -140 6870
rect -90 6830 100 6870
rect 150 6830 340 6870
rect 390 6830 580 6870
rect 3140 6830 3330 6870
rect 3380 6830 3570 6870
rect 3620 6830 3810 6870
rect 3860 6830 4050 6870
rect 740 6320 780 6360
rect 880 6320 920 6360
rect 1460 6320 1500 6360
rect 2220 6320 2260 6360
rect 2940 6320 2980 6360
rect 4320 6400 4360 6440
rect -330 5840 -140 5880
rect 1840 5790 1880 5830
rect 3860 5840 4050 5880
rect 1590 5700 1650 5750
rect 2070 5700 2130 5750
rect 870 5620 930 5670
rect 2790 5620 2850 5670
rect 760 5200 800 5240
rect 1830 5260 1890 5310
rect 1480 5200 1520 5240
rect 2200 5200 2240 5240
rect 2920 5230 2960 5270
rect -330 4770 -140 4810
rect 1840 4730 1880 4770
rect 3860 4770 4050 4810
<< locali >>
rect 3980 10000 4060 10020
rect 3980 9960 4000 10000
rect 4040 9990 4060 10000
rect 4040 9960 4260 9990
rect 3980 9940 4260 9960
rect 850 9900 2870 9940
rect 850 9830 950 9900
rect -450 9790 950 9830
rect -450 6660 -410 9790
rect -350 9620 -250 9640
rect -350 9380 -330 9620
rect -270 9380 -250 9620
rect -350 9320 -250 9380
rect -110 9620 -10 9640
rect -110 9380 -90 9620
rect -30 9380 -10 9620
rect -110 9320 -10 9380
rect 130 9620 230 9640
rect 130 9380 150 9620
rect 210 9380 230 9620
rect 130 9320 230 9380
rect 370 9620 470 9640
rect 370 9380 390 9620
rect 450 9380 470 9620
rect 370 9320 470 9380
rect 610 9620 710 9640
rect 610 9380 630 9620
rect 690 9380 710 9620
rect 610 9320 710 9380
rect 850 9620 950 9790
rect 850 9380 870 9620
rect 930 9380 950 9620
rect 850 9360 950 9380
rect 1090 9820 2630 9860
rect 1090 9620 1190 9820
rect 1230 9750 1310 9780
rect 1230 9710 1250 9750
rect 1290 9710 1310 9750
rect 1230 9680 1310 9710
rect 1090 9380 1110 9620
rect 1170 9380 1190 9620
rect 1090 9360 1190 9380
rect 1330 9620 1430 9640
rect 1330 9380 1350 9620
rect 1410 9380 1430 9620
rect -350 9300 840 9320
rect -350 9260 -330 9300
rect -140 9260 -90 9300
rect 100 9260 150 9300
rect 340 9260 390 9300
rect 580 9260 630 9300
rect 820 9260 840 9300
rect -350 9240 840 9260
rect 1330 9270 1430 9380
rect 1570 9620 1670 9820
rect 1570 9380 1590 9620
rect 1650 9380 1670 9620
rect 1570 9360 1670 9380
rect 1810 9620 1910 9640
rect 1810 9380 1830 9620
rect 1890 9380 1910 9620
rect 1810 9360 1910 9380
rect 2050 9620 2150 9820
rect 2410 9750 2490 9780
rect 2410 9710 2430 9750
rect 2470 9710 2490 9750
rect 2410 9680 2490 9710
rect 2050 9380 2070 9620
rect 2130 9380 2150 9620
rect 2050 9360 2150 9380
rect 2290 9620 2390 9640
rect 2290 9380 2310 9620
rect 2370 9380 2390 9620
rect 2290 9270 2390 9380
rect 2530 9620 2630 9820
rect 2530 9380 2550 9620
rect 2610 9380 2630 9620
rect 2530 9360 2630 9380
rect 2770 9620 2870 9900
rect 2770 9380 2790 9620
rect 2850 9380 2870 9620
rect 2770 9360 2870 9380
rect 3010 9620 3110 9640
rect 3010 9380 3030 9620
rect 3090 9380 3110 9620
rect 3010 9320 3110 9380
rect 3250 9620 3350 9640
rect 3250 9380 3270 9620
rect 3330 9380 3350 9620
rect 3250 9320 3350 9380
rect 3490 9620 3590 9640
rect 3490 9380 3510 9620
rect 3570 9380 3590 9620
rect 3490 9320 3590 9380
rect 3730 9620 3830 9640
rect 3730 9380 3750 9620
rect 3810 9380 3830 9620
rect 3730 9320 3830 9380
rect 3970 9620 4070 9640
rect 3970 9380 3990 9620
rect 4050 9380 4070 9620
rect 3970 9320 4070 9380
rect 1330 9230 2390 9270
rect 2880 9300 4070 9320
rect 2880 9260 2900 9300
rect 3090 9260 3140 9300
rect 3330 9260 3380 9300
rect 3570 9260 3620 9300
rect 3810 9260 3860 9300
rect 4050 9260 4070 9300
rect 2880 9240 4070 9260
rect 710 9190 810 9200
rect 340 9150 440 9170
rect 340 9090 360 9150
rect 420 9090 440 9150
rect 710 9130 730 9190
rect 790 9130 810 9190
rect 710 9110 810 9130
rect 1540 9190 1630 9230
rect 1540 9140 1560 9190
rect 1610 9140 1630 9190
rect 2930 9190 3030 9200
rect 1540 9120 1630 9140
rect 1820 9160 1900 9180
rect 1820 9120 1840 9160
rect 1880 9140 1900 9160
rect 1880 9120 2470 9140
rect 1820 9100 2470 9120
rect 2930 9130 2950 9190
rect 3010 9130 3030 9190
rect 2930 9110 3030 9130
rect 3450 9180 3550 9200
rect 3450 9120 3470 9180
rect 3530 9120 3550 9180
rect 3450 9100 3550 9120
rect 340 9070 440 9090
rect 2430 9060 2470 9100
rect 4040 9080 4120 9100
rect 4040 9060 4060 9080
rect 1330 9020 2390 9060
rect 2430 9040 4060 9060
rect 4100 9040 4120 9080
rect 2430 9020 4120 9040
rect -350 8960 -250 8980
rect -350 8720 -330 8960
rect -270 8720 -250 8960
rect -350 8660 -250 8720
rect -110 8960 -10 8980
rect -110 8720 -90 8960
rect -30 8720 -10 8960
rect -110 8660 -10 8720
rect 130 8960 230 8980
rect 130 8720 150 8960
rect 210 8720 230 8960
rect 130 8660 230 8720
rect 370 8960 470 8980
rect 370 8720 390 8960
rect 450 8720 470 8960
rect 370 8660 470 8720
rect 610 8960 710 8980
rect 610 8720 630 8960
rect 690 8720 710 8960
rect 610 8660 710 8720
rect 850 8960 950 8980
rect 850 8720 870 8960
rect 930 8720 950 8960
rect 850 8700 950 8720
rect -350 8640 840 8660
rect -350 8600 -330 8640
rect -140 8600 -90 8640
rect 100 8600 150 8640
rect 340 8600 390 8640
rect 580 8600 630 8640
rect 820 8600 840 8640
rect -350 8580 840 8600
rect 910 8470 950 8700
rect 1090 8960 1190 8980
rect 1090 8720 1110 8960
rect 1170 8720 1190 8960
rect 1090 8550 1190 8720
rect 1330 8960 1430 9020
rect 1330 8720 1350 8960
rect 1410 8720 1430 8960
rect 1330 8700 1430 8720
rect 1570 8960 1670 8980
rect 1570 8720 1590 8960
rect 1650 8720 1670 8960
rect 1450 8650 1530 8670
rect 1450 8610 1470 8650
rect 1510 8610 1530 8650
rect 1450 8590 1530 8610
rect 1570 8550 1670 8720
rect 1810 8960 1910 8980
rect 1810 8720 1830 8960
rect 1890 8720 1910 8960
rect 1810 8700 1910 8720
rect 2050 8960 2150 8980
rect 2050 8720 2070 8960
rect 2130 8720 2150 8960
rect 2050 8550 2150 8720
rect 2290 8960 2390 9020
rect 2290 8720 2310 8960
rect 2370 8720 2390 8960
rect 2290 8700 2390 8720
rect 2530 8960 2630 8980
rect 2530 8720 2550 8960
rect 2610 8720 2630 8960
rect 2190 8650 2270 8670
rect 2190 8610 2210 8650
rect 2250 8610 2270 8650
rect 2190 8590 2270 8610
rect 2320 8640 2380 8700
rect 2320 8600 2330 8640
rect 2370 8600 2380 8640
rect 2320 8590 2380 8600
rect 2530 8550 2630 8720
rect 1090 8510 2630 8550
rect 2770 8960 2870 8980
rect 2770 8720 2790 8960
rect 2850 8720 2870 8960
rect 2770 8700 2870 8720
rect 3010 8960 3110 8980
rect 3010 8720 3030 8960
rect 3090 8720 3110 8960
rect 2770 8470 2810 8700
rect 3010 8660 3110 8720
rect 3250 8960 3350 8980
rect 3250 8720 3270 8960
rect 3330 8720 3350 8960
rect 3250 8660 3350 8720
rect 3490 8960 3590 8980
rect 3490 8720 3510 8960
rect 3570 8720 3590 8960
rect 3490 8660 3590 8720
rect 3730 8960 3830 8980
rect 3730 8720 3750 8960
rect 3810 8720 3830 8960
rect 3730 8660 3830 8720
rect 3970 8960 4070 8980
rect 3970 8720 3990 8960
rect 4050 8720 4070 8960
rect 3970 8660 4070 8720
rect 2880 8640 4070 8660
rect 2880 8600 2900 8640
rect 3090 8600 3140 8640
rect 3330 8600 3380 8640
rect 3570 8600 3620 8640
rect 3810 8600 3860 8640
rect 4050 8600 4070 8640
rect 2880 8580 4070 8600
rect 910 8430 2810 8470
rect 910 8390 950 8430
rect 2770 8390 2810 8430
rect 910 8350 4160 8390
rect 910 8100 950 8350
rect -350 8070 -250 8090
rect -350 7830 -330 8070
rect -270 7830 -250 8070
rect -350 7770 -250 7830
rect -110 8070 -10 8090
rect -110 7830 -90 8070
rect -30 7830 -10 8070
rect -110 7770 -10 7830
rect 130 8070 230 8090
rect 130 7830 150 8070
rect 210 7830 230 8070
rect 130 7770 230 7830
rect 370 8070 470 8090
rect 370 7830 390 8070
rect 450 7830 470 8070
rect 370 7770 470 7830
rect 610 8070 710 8090
rect 610 7830 630 8070
rect 690 7830 710 8070
rect 610 7810 710 7830
rect 850 8070 950 8100
rect 1570 8300 2380 8310
rect 1570 8270 2330 8300
rect 850 7830 870 8070
rect 930 7830 950 8070
rect 850 7810 950 7830
rect 1090 8070 1190 8090
rect 1090 7830 1110 8070
rect 1170 7830 1190 8070
rect 1090 7770 1190 7830
rect 1330 8070 1430 8090
rect 1330 7830 1350 8070
rect 1410 7830 1430 8070
rect 1330 7770 1430 7830
rect 1570 8070 1670 8270
rect 2050 8260 2330 8270
rect 2370 8260 2380 8300
rect 2050 8250 2380 8260
rect 1570 7830 1590 8070
rect 1650 7830 1670 8070
rect 1570 7810 1670 7830
rect 1810 8070 1910 8090
rect 1810 7830 1830 8070
rect 1890 7830 1910 8070
rect 1810 7810 1910 7830
rect 2050 8070 2150 8250
rect 2770 8100 2810 8350
rect 2050 7830 2070 8070
rect 2130 7830 2150 8070
rect 2050 7810 2150 7830
rect 2290 8070 2390 8090
rect 2290 7830 2310 8070
rect 2370 7830 2390 8070
rect -350 7750 600 7770
rect -350 7710 -330 7750
rect -140 7710 -90 7750
rect 100 7710 150 7750
rect 340 7710 390 7750
rect 580 7710 600 7750
rect -350 7690 600 7710
rect 960 7750 1190 7770
rect 960 7710 980 7750
rect 1060 7710 1190 7750
rect 960 7690 1190 7710
rect 1240 7750 1430 7770
rect 1240 7710 1260 7750
rect 1300 7730 1430 7750
rect 1680 7750 1800 7770
rect 1300 7710 1320 7730
rect 1240 7690 1320 7710
rect 1680 7710 1700 7750
rect 1780 7710 1800 7750
rect 1680 7690 1800 7710
rect 730 7670 830 7690
rect 730 7600 750 7670
rect 810 7600 830 7670
rect 730 7580 830 7600
rect 960 7530 1080 7690
rect 1680 7530 1780 7690
rect 1840 7650 1880 7810
rect 2290 7770 2390 7830
rect 2530 8070 2630 8090
rect 2530 7830 2550 8070
rect 2610 7830 2630 8070
rect 2530 7770 2630 7830
rect 2770 8070 2870 8100
rect 2770 7830 2790 8070
rect 2850 7830 2870 8070
rect 2770 7810 2870 7830
rect 3010 8070 3110 8090
rect 3010 7830 3030 8070
rect 3090 7830 3110 8070
rect 3010 7810 3110 7830
rect 3250 8070 3350 8090
rect 3250 7830 3270 8070
rect 3330 7830 3350 8070
rect 3250 7770 3350 7830
rect 3490 8070 3590 8090
rect 3490 7830 3510 8070
rect 3570 7830 3590 8070
rect 3490 7770 3590 7830
rect 3730 8070 3830 8090
rect 3730 7830 3750 8070
rect 3810 7830 3830 8070
rect 3730 7770 3830 7830
rect 3970 8070 4070 8090
rect 3970 7830 3990 8070
rect 4050 7830 4070 8070
rect 3970 7770 4070 7830
rect 1920 7750 2040 7770
rect 1920 7710 1940 7750
rect 2020 7710 2040 7750
rect 2290 7750 2480 7770
rect 2290 7730 2420 7750
rect 1920 7690 2040 7710
rect 2400 7710 2420 7730
rect 2460 7710 2480 7750
rect 2400 7690 2480 7710
rect 2530 7750 2760 7770
rect 2530 7710 2660 7750
rect 2740 7710 2760 7750
rect 2530 7690 2760 7710
rect 3120 7750 4070 7770
rect 3120 7710 3140 7750
rect 3330 7710 3380 7750
rect 3570 7710 3620 7750
rect 3810 7710 3860 7750
rect 4050 7710 4070 7750
rect 3120 7690 4070 7710
rect 1820 7630 1900 7650
rect 1820 7590 1840 7630
rect 1880 7590 1900 7630
rect 1820 7570 1900 7590
rect 1940 7530 2040 7690
rect 2640 7530 2760 7690
rect 2890 7650 2990 7670
rect 2890 7580 2910 7650
rect 2970 7580 2990 7650
rect 4120 7590 4160 8350
rect 2890 7560 2990 7580
rect 340 7510 440 7530
rect 340 7440 360 7510
rect 420 7440 440 7510
rect 340 7420 440 7440
rect 960 7490 2760 7530
rect 3900 7550 4160 7590
rect 960 7330 1080 7490
rect 1560 7370 1640 7400
rect 1560 7330 1580 7370
rect 1620 7330 1640 7370
rect 960 7310 1190 7330
rect 960 7270 980 7310
rect 1060 7270 1190 7310
rect 960 7250 1190 7270
rect 1240 7310 1320 7330
rect 1240 7270 1260 7310
rect 1300 7290 1320 7310
rect 1560 7300 1640 7330
rect 1300 7270 1430 7290
rect 1240 7250 1430 7270
rect -350 7190 -250 7210
rect -350 6950 -330 7190
rect -270 6950 -250 7190
rect -350 6890 -250 6950
rect -110 7190 -10 7210
rect -110 6950 -90 7190
rect -30 6950 -10 7190
rect -110 6890 -10 6950
rect 130 7190 230 7210
rect 130 6950 150 7190
rect 210 6950 230 7190
rect 130 6890 230 6950
rect 370 7190 470 7210
rect 370 6950 390 7190
rect 450 6950 470 7190
rect 370 6890 470 6950
rect 610 7190 710 7210
rect 610 6950 630 7190
rect 690 6950 710 7190
rect 610 6930 710 6950
rect 850 7190 950 7210
rect 850 6950 870 7190
rect 930 6950 950 7190
rect -350 6870 600 6890
rect -350 6830 -330 6870
rect -140 6830 -90 6870
rect 100 6830 150 6870
rect 340 6830 390 6870
rect 580 6830 600 6870
rect -350 6810 600 6830
rect 850 6660 950 6950
rect 1090 7190 1190 7250
rect 1090 6950 1110 7190
rect 1170 6950 1190 7190
rect 1090 6930 1190 6950
rect 1330 7190 1430 7250
rect 1330 6950 1350 7190
rect 1410 6950 1430 7190
rect 1330 6930 1430 6950
rect 1570 7210 1640 7300
rect 1680 7330 1780 7490
rect 1820 7430 1900 7450
rect 1820 7390 1840 7430
rect 1880 7390 1900 7430
rect 1820 7370 1900 7390
rect 1680 7310 1800 7330
rect 1680 7270 1700 7310
rect 1780 7270 1800 7310
rect 1680 7250 1800 7270
rect 1840 7210 1880 7370
rect 1940 7330 2040 7490
rect 2640 7330 2760 7490
rect 3360 7490 3460 7510
rect 3360 7420 3380 7490
rect 3440 7420 3460 7490
rect 3360 7400 3460 7420
rect 3900 7390 3950 7550
rect 4220 7510 4260 9940
rect 3990 7490 4260 7510
rect 3990 7450 4010 7490
rect 4050 7470 4260 7490
rect 4050 7450 4070 7470
rect 3990 7430 4070 7450
rect 3900 7350 4160 7390
rect 1920 7310 2040 7330
rect 1920 7270 1940 7310
rect 2020 7270 2040 7310
rect 2400 7310 2480 7330
rect 2400 7290 2420 7310
rect 1920 7250 2040 7270
rect 2290 7270 2420 7290
rect 2460 7270 2480 7310
rect 2290 7250 2480 7270
rect 2530 7310 2760 7330
rect 2530 7270 2660 7310
rect 2740 7270 2760 7310
rect 2530 7250 2760 7270
rect 1570 7190 1670 7210
rect 1570 6950 1590 7190
rect 1650 6950 1670 7190
rect 1570 6740 1670 6950
rect 1810 7190 1910 7210
rect 1810 6950 1830 7190
rect 1890 6950 1910 7190
rect 1810 6930 1910 6950
rect 2050 7190 2150 7210
rect 2050 6950 2070 7190
rect 2130 6950 2150 7190
rect 2050 6740 2150 6950
rect 2290 7190 2390 7250
rect 2290 6950 2310 7190
rect 2370 6950 2390 7190
rect 2290 6930 2390 6950
rect 2530 7190 2630 7250
rect 2530 6950 2550 7190
rect 2610 6950 2630 7190
rect 2530 6930 2630 6950
rect 2770 7190 2870 7210
rect 2770 6950 2790 7190
rect 2850 6950 2870 7190
rect 1570 6700 2150 6740
rect 2770 6660 2870 6950
rect 3010 7190 3110 7210
rect 3010 6950 3030 7190
rect 3090 6950 3110 7190
rect 3010 6930 3110 6950
rect 3250 7190 3350 7210
rect 3250 6950 3270 7190
rect 3330 6950 3350 7190
rect 3250 6890 3350 6950
rect 3490 7190 3590 7210
rect 3490 6950 3510 7190
rect 3570 6950 3590 7190
rect 3490 6890 3590 6950
rect 3730 7190 3830 7210
rect 3730 6950 3750 7190
rect 3810 6950 3830 7190
rect 3730 6890 3830 6950
rect 3970 7190 4070 7210
rect 3970 6950 3990 7190
rect 4050 6950 4070 7190
rect 3970 6890 4070 6950
rect 3120 6870 4070 6890
rect 3120 6830 3140 6870
rect 3330 6830 3380 6870
rect 3570 6830 3620 6870
rect 3810 6830 3860 6870
rect 4050 6830 4070 6870
rect 3120 6810 4070 6830
rect -450 6640 2870 6660
rect -450 6620 1840 6640
rect 1820 6600 1840 6620
rect 1880 6620 2870 6640
rect 1880 6600 1900 6620
rect 1820 6580 1900 6600
rect 4120 6580 4160 7350
rect 2060 6560 4160 6580
rect 2060 6520 2080 6560
rect 2120 6520 4160 6560
rect 2060 6500 4160 6520
rect 4220 6460 4260 7470
rect 130 6420 3590 6460
rect 4220 6440 4380 6460
rect 4220 6420 4320 6440
rect -350 6200 -250 6220
rect -350 5960 -330 6200
rect -270 5960 -250 6200
rect -350 5900 -250 5960
rect -110 6200 -10 6220
rect -110 5960 -90 6200
rect -30 5960 -10 6200
rect -110 5940 -10 5960
rect 130 6200 230 6420
rect 610 6230 650 6420
rect 720 6360 800 6380
rect 720 6320 740 6360
rect 780 6320 800 6360
rect 720 6300 800 6320
rect 860 6360 940 6380
rect 860 6320 880 6360
rect 920 6320 940 6360
rect 860 6300 940 6320
rect 130 5960 150 6200
rect 210 5960 230 6200
rect 130 5940 230 5960
rect 370 6200 470 6220
rect 370 5960 390 6200
rect 450 5960 470 6200
rect 370 5940 470 5960
rect 610 6200 710 6230
rect 610 5960 630 6200
rect 690 5960 710 6200
rect 610 5940 710 5960
rect 850 6200 950 6300
rect 850 5960 870 6200
rect 930 5960 950 6200
rect -350 5880 -120 5900
rect -350 5840 -330 5880
rect -140 5840 -120 5880
rect -350 5820 -120 5840
rect 480 5740 700 5760
rect 480 5560 500 5740
rect 680 5560 700 5740
rect 850 5670 950 5960
rect 1090 6200 1190 6420
rect 1440 6360 1520 6380
rect 1440 6320 1460 6360
rect 1500 6320 1520 6360
rect 1440 6300 1520 6320
rect 2200 6360 2280 6380
rect 2200 6320 2220 6360
rect 2260 6320 2280 6360
rect 2200 6300 2280 6320
rect 1090 5960 1110 6200
rect 1170 5960 1190 6200
rect 1090 5940 1190 5960
rect 1330 6200 1430 6220
rect 1330 5960 1350 6200
rect 1410 5960 1430 6200
rect 1330 5940 1430 5960
rect 1570 6200 1670 6220
rect 1570 5960 1590 6200
rect 1650 5960 1670 6200
rect 1570 5750 1670 5960
rect 1570 5700 1590 5750
rect 1650 5700 1670 5750
rect 1570 5680 1670 5700
rect 1810 6200 1910 6220
rect 1810 5960 1830 6200
rect 1890 5960 1910 6200
rect 1810 5830 1910 5960
rect 1810 5790 1840 5830
rect 1880 5790 1910 5830
rect 850 5620 870 5670
rect 930 5620 950 5670
rect 850 5600 950 5620
rect 480 5540 700 5560
rect 1810 5510 1910 5790
rect 2050 6200 2150 6220
rect 2050 5960 2070 6200
rect 2130 5960 2150 6200
rect 2050 5750 2150 5960
rect 2290 6200 2390 6220
rect 2290 5960 2310 6200
rect 2370 5960 2390 6200
rect 2290 5940 2390 5960
rect 2530 6200 2630 6420
rect 2920 6360 3000 6380
rect 2920 6320 2940 6360
rect 2980 6320 3000 6360
rect 2920 6300 3000 6320
rect 3070 6230 3110 6420
rect 2530 5960 2550 6200
rect 2610 5960 2630 6200
rect 2530 5940 2630 5960
rect 2770 6200 2870 6220
rect 2770 5960 2790 6200
rect 2850 5960 2870 6200
rect 2050 5700 2070 5750
rect 2130 5700 2150 5750
rect 2050 5680 2150 5700
rect 2770 5670 2870 5960
rect 3010 6200 3110 6230
rect 3010 5960 3030 6200
rect 3090 5960 3110 6200
rect 3010 5940 3110 5960
rect 3250 6200 3350 6220
rect 3250 5960 3270 6200
rect 3330 5960 3350 6200
rect 3250 5940 3350 5960
rect 3490 6200 3590 6420
rect 4300 6400 4320 6420
rect 4360 6400 4380 6440
rect 4300 6380 4380 6400
rect 5240 6420 5330 6440
rect 5240 6370 5260 6420
rect 5310 6370 5330 6420
rect 3490 5960 3510 6200
rect 3570 5960 3590 6200
rect 3490 5940 3590 5960
rect 3730 6200 3830 6220
rect 3730 5960 3750 6200
rect 3810 5960 3830 6200
rect 3730 5940 3830 5960
rect 3970 6200 4070 6220
rect 3970 5960 3990 6200
rect 4050 5960 4070 6200
rect 3970 5900 4070 5960
rect 3840 5880 4070 5900
rect 3840 5840 3860 5880
rect 4050 5840 4070 5880
rect 3840 5820 4070 5840
rect 5240 5820 5330 6370
rect 5170 5770 5420 5820
rect 2770 5620 2790 5670
rect 2850 5620 2870 5670
rect 2770 5600 2870 5620
rect 3040 5740 3260 5760
rect 3040 5560 3060 5740
rect 3240 5560 3260 5740
rect 3040 5540 3260 5560
rect 910 5460 1130 5480
rect 910 5280 930 5460
rect 1110 5280 1130 5460
rect 910 5260 1130 5280
rect 1330 5470 2390 5510
rect 740 5240 820 5260
rect 740 5200 760 5240
rect 800 5200 820 5240
rect 740 5180 820 5200
rect 1330 5160 1370 5470
rect 1630 5390 1840 5410
rect 1880 5390 2090 5410
rect 1630 5370 2090 5390
rect 1460 5240 1540 5260
rect 1460 5200 1480 5240
rect 1520 5200 1540 5240
rect 1460 5180 1540 5200
rect 1630 5160 1670 5370
rect -350 5130 -250 5150
rect -350 4890 -330 5130
rect -270 4890 -250 5130
rect -350 4830 -250 4890
rect -110 5130 -10 5150
rect -110 4890 -90 5130
rect -30 4890 -10 5130
rect -110 4870 -10 4890
rect 130 5130 230 5150
rect 130 4890 150 5130
rect 210 4890 230 5130
rect -350 4810 -120 4830
rect -350 4770 -330 4810
rect -140 4770 -120 4810
rect -350 4750 -120 4770
rect 130 4670 230 4890
rect 370 5130 470 5150
rect 370 4890 390 5130
rect 450 4890 470 5130
rect 370 4870 470 4890
rect 610 5130 710 5150
rect 610 4890 630 5130
rect 690 4890 710 5130
rect 610 4670 710 4890
rect 850 5130 950 5150
rect 850 4890 870 5130
rect 930 4890 950 5130
rect 850 4870 950 4890
rect 1090 5130 1190 5150
rect 1090 4890 1110 5130
rect 1170 4890 1190 5130
rect 1090 4670 1190 4890
rect 1330 5130 1430 5160
rect 1330 4890 1350 5130
rect 1410 4890 1430 5130
rect 1330 4870 1430 4890
rect 1570 5130 1670 5160
rect 1570 4890 1590 5130
rect 1650 4890 1670 5130
rect 1570 4870 1670 4890
rect 1810 5310 1910 5330
rect 1810 5260 1830 5310
rect 1890 5260 1910 5310
rect 1810 5130 1910 5260
rect 1810 4890 1830 5130
rect 1890 4890 1910 5130
rect 1810 4870 1910 4890
rect 2050 5160 2090 5370
rect 2180 5240 2260 5260
rect 2180 5200 2200 5240
rect 2240 5200 2260 5240
rect 2180 5180 2260 5200
rect 2350 5160 2390 5470
rect 2590 5460 2810 5480
rect 2590 5280 2610 5460
rect 2790 5280 2810 5460
rect 2590 5260 2810 5280
rect 2900 5270 2980 5290
rect 2900 5230 2920 5270
rect 2960 5230 2980 5270
rect 2900 5210 2980 5230
rect 2050 5130 2150 5160
rect 2050 4890 2070 5130
rect 2130 4890 2150 5130
rect 2050 4870 2150 4890
rect 2290 5130 2390 5160
rect 2290 4890 2310 5130
rect 2370 4890 2390 5130
rect 2290 4870 2390 4890
rect 2530 5130 2630 5150
rect 2530 4890 2550 5130
rect 2610 4890 2630 5130
rect 1820 4770 1900 4870
rect 1820 4730 1840 4770
rect 1880 4730 1900 4770
rect 1820 4710 1900 4730
rect 2530 4670 2630 4890
rect 2770 5130 2870 5150
rect 2770 4890 2790 5130
rect 2850 4890 2870 5130
rect 2770 4870 2870 4890
rect 3010 5130 3110 5150
rect 3010 4890 3030 5130
rect 3090 4890 3110 5130
rect 3010 4670 3110 4890
rect 3250 5130 3350 5150
rect 3250 4890 3270 5130
rect 3330 4890 3350 5130
rect 3250 4870 3350 4890
rect 3490 5130 3590 5150
rect 3490 4890 3510 5130
rect 3570 4890 3590 5130
rect 3490 4670 3590 4890
rect 3730 5130 3830 5150
rect 3730 4890 3750 5130
rect 3810 4890 3830 5130
rect 3730 4870 3830 4890
rect 3970 5130 4070 5150
rect 3970 4890 3990 5130
rect 4050 4890 4070 5130
rect 3970 4830 4070 4890
rect 3840 4810 4070 4830
rect 3840 4770 3860 4810
rect 4050 4770 4070 4810
rect 3840 4750 4070 4770
rect 130 4630 3590 4670
<< viali >>
rect 4000 9960 4040 10000
rect -330 9380 -270 9620
rect -90 9380 -30 9620
rect 150 9380 210 9620
rect 390 9380 450 9620
rect 630 9380 690 9620
rect 1250 9710 1290 9750
rect 1830 9380 1890 9620
rect 2430 9710 2470 9750
rect 3030 9380 3090 9620
rect 3270 9380 3330 9620
rect 3510 9380 3570 9620
rect 3750 9380 3810 9620
rect 3990 9380 4050 9620
rect 360 9090 420 9150
rect 730 9130 790 9190
rect 1560 9140 1610 9190
rect 2950 9130 3010 9190
rect 3470 9120 3530 9180
rect -330 8720 -270 8960
rect -90 8720 -30 8960
rect 150 8720 210 8960
rect 390 8720 450 8960
rect 1470 8610 1510 8650
rect 1830 8720 1890 8960
rect 2210 8610 2250 8650
rect 2330 8600 2370 8640
rect 3270 8720 3330 8960
rect 3510 8720 3570 8960
rect 3750 8720 3810 8960
rect 3990 8720 4050 8960
rect -330 7830 -270 8070
rect -90 7830 -30 8070
rect 150 7830 210 8070
rect 390 7830 450 8070
rect 630 7830 690 8070
rect 1350 7830 1410 8070
rect 2330 8260 2370 8300
rect 2310 7830 2370 8070
rect 750 7600 810 7670
rect 3030 7830 3090 8070
rect 3270 7830 3330 8070
rect 3510 7830 3570 8070
rect 3750 7830 3810 8070
rect 3990 7830 4050 8070
rect 2910 7580 2970 7650
rect 360 7440 420 7510
rect 1580 7330 1620 7370
rect -330 6950 -270 7190
rect -90 6950 -30 7190
rect 150 6950 210 7190
rect 390 6950 450 7190
rect 630 6950 690 7190
rect 1350 6950 1410 7190
rect 3380 7420 3440 7490
rect 2310 6950 2370 7190
rect 3030 6950 3090 7190
rect 3270 6950 3330 7190
rect 3510 6950 3570 7190
rect 3750 6950 3810 7190
rect 3990 6950 4050 7190
rect 1840 6600 1880 6640
rect 2080 6520 2120 6560
rect -330 5960 -270 6200
rect -90 5960 -30 6200
rect 740 6320 780 6360
rect 390 5960 450 6200
rect 500 5560 680 5740
rect 1460 6320 1500 6360
rect 2220 6320 2260 6360
rect 1350 5960 1410 6200
rect 2310 5960 2370 6200
rect 2940 6320 2980 6360
rect 2070 5700 2130 5750
rect 3270 5960 3330 6200
rect 5260 6370 5310 6420
rect 3750 5960 3810 6200
rect 3990 5960 4050 6200
rect 3060 5560 3240 5740
rect 930 5280 1110 5460
rect 760 5200 800 5240
rect 1840 5390 1880 5430
rect 1480 5200 1520 5240
rect -330 4890 -270 5130
rect -90 4890 -30 5130
rect 390 4890 450 5130
rect 870 4890 930 5130
rect 2200 5200 2240 5240
rect 2610 5280 2790 5460
rect 2920 5230 2960 5270
rect 2790 4890 2850 5130
rect 3270 4890 3330 5130
rect 3750 4890 3810 5130
rect 3990 4890 4050 5130
<< metal1 >>
rect 3980 10010 4060 10020
rect 3980 9950 3990 10010
rect 4050 9950 4060 10010
rect 3980 9940 4060 9950
rect 1210 9760 1310 9780
rect 1210 9700 1240 9760
rect 1300 9700 1310 9760
rect 1210 9660 1310 9700
rect 2410 9760 2510 9780
rect 2410 9700 2420 9760
rect 2480 9700 2510 9760
rect 2410 9660 2510 9700
rect -350 9620 -250 9640
rect -350 9380 -330 9620
rect -270 9380 -250 9620
rect -350 9360 -250 9380
rect -110 9620 -10 9640
rect -110 9380 -90 9620
rect -30 9380 -10 9620
rect -110 9360 -10 9380
rect 130 9620 230 9640
rect 130 9380 150 9620
rect 210 9380 230 9620
rect 130 9360 230 9380
rect 370 9620 470 9640
rect 370 9380 390 9620
rect 450 9380 470 9620
rect 370 9360 470 9380
rect 610 9620 710 9640
rect 610 9380 630 9620
rect 690 9380 710 9620
rect 610 9360 710 9380
rect 840 9360 1190 9640
rect 1810 9620 1910 9640
rect 1810 9380 1830 9620
rect 1890 9380 1910 9620
rect 1810 9360 1910 9380
rect 2530 9360 2880 9640
rect 3010 9620 3110 9640
rect 3010 9380 3030 9620
rect 3090 9380 3110 9620
rect 3010 9360 3110 9380
rect 3250 9620 3350 9640
rect 3250 9380 3270 9620
rect 3330 9380 3350 9620
rect 3250 9360 3350 9380
rect 3490 9620 3590 9640
rect 3490 9380 3510 9620
rect 3570 9380 3590 9620
rect 3490 9360 3590 9380
rect 3730 9620 3830 9640
rect 3730 9380 3750 9620
rect 3810 9380 3830 9620
rect 3730 9360 3830 9380
rect 3970 9620 4070 9640
rect 3970 9380 3990 9620
rect 4050 9380 4070 9620
rect 3970 9360 4070 9380
rect 700 9190 820 9210
rect 330 9150 450 9180
rect 330 9090 360 9150
rect 420 9090 450 9150
rect 700 9130 730 9190
rect 790 9130 820 9190
rect 700 9100 820 9130
rect 330 8980 450 9090
rect 1090 8980 1190 9360
rect 1540 9190 1630 9210
rect 1540 9140 1560 9190
rect 1610 9140 1630 9190
rect 1540 9090 1630 9140
rect 1540 9060 1700 9090
rect -510 8960 1560 8980
rect -510 8720 -330 8960
rect -270 8720 -90 8960
rect -30 8720 150 8960
rect 210 8720 390 8960
rect 450 8720 1560 8960
rect -510 8700 1560 8720
rect -510 7540 -410 8700
rect 1440 8650 1560 8700
rect 1440 8610 1470 8650
rect 1510 8610 1560 8650
rect 1440 8590 1560 8610
rect -350 8070 -250 8090
rect -350 7830 -330 8070
rect -270 7830 -250 8070
rect -350 7810 -250 7830
rect -110 8070 -10 8090
rect -110 7830 -90 8070
rect -30 7830 -10 8070
rect -110 7810 -10 7830
rect 130 8070 230 8090
rect 130 7830 150 8070
rect 210 7830 230 8070
rect 130 7810 230 7830
rect 370 8070 470 8090
rect 370 7830 390 8070
rect 450 7830 470 8070
rect 370 7810 470 7830
rect 610 8070 710 8080
rect 610 7830 630 8070
rect 690 7830 710 8070
rect 610 7810 710 7830
rect 1330 8070 1430 8090
rect 1330 7830 1350 8070
rect 1410 7830 1430 8070
rect 1330 7810 1430 7830
rect 730 7670 830 7690
rect 730 7600 750 7670
rect 810 7600 830 7670
rect 730 7580 830 7600
rect 1600 7550 1700 9060
rect 2530 8980 2630 9360
rect 2920 9190 3040 9210
rect 2920 9130 2950 9190
rect 3010 9130 3040 9190
rect 2920 9100 3040 9130
rect 3440 9180 3560 9210
rect 3440 9120 3470 9180
rect 3530 9120 3560 9180
rect 3440 8980 3560 9120
rect 1810 8960 4220 8980
rect 1810 8720 1830 8960
rect 1890 8720 3270 8960
rect 3330 8720 3510 8960
rect 3570 8720 3750 8960
rect 3810 8720 3990 8960
rect 4050 8720 4220 8960
rect 1810 8700 4220 8720
rect 2160 8650 2280 8700
rect 2160 8610 2210 8650
rect 2250 8610 2280 8650
rect 2160 8590 2280 8610
rect 2310 8640 2390 8660
rect 2310 8600 2330 8640
rect 2370 8600 2390 8640
rect 2310 8300 2390 8600
rect 2310 8260 2330 8300
rect 2370 8260 2390 8300
rect 2310 8240 2390 8260
rect 2290 8070 2390 8090
rect 2290 7830 2310 8070
rect 2370 7830 2390 8070
rect 2290 7810 2390 7830
rect 3010 8070 3110 8090
rect 3010 7830 3030 8070
rect 3090 7830 3110 8070
rect 3010 7810 3110 7830
rect 3250 8070 3350 8090
rect 3250 7830 3270 8070
rect 3330 7830 3350 8070
rect 3250 7810 3350 7830
rect 3490 8070 3590 8090
rect 3490 7830 3510 8070
rect 3570 7830 3590 8070
rect 3490 7810 3590 7830
rect 3730 8070 3830 8090
rect 3730 7830 3750 8070
rect 3810 7830 3830 8070
rect 3730 7810 3830 7830
rect 3970 8070 4070 8090
rect 3970 7830 3990 8070
rect 4050 7830 4070 8070
rect 3970 7810 4070 7830
rect 2890 7650 2990 7670
rect 2890 7580 2910 7650
rect 2970 7580 2990 7650
rect 2890 7560 2990 7580
rect -510 7510 450 7540
rect -510 7440 360 7510
rect 420 7440 450 7510
rect -510 7410 450 7440
rect 330 7210 450 7410
rect 1560 7470 1700 7550
rect 4120 7520 4220 8700
rect 3350 7490 4220 7520
rect 1560 7370 1640 7470
rect 1560 7330 1580 7370
rect 1620 7330 1640 7370
rect 1560 7300 1640 7330
rect 3350 7420 3380 7490
rect 3440 7420 4220 7490
rect 3350 7390 4220 7420
rect 3350 7210 3470 7390
rect -360 7190 1430 7210
rect -360 6950 -330 7190
rect -270 6950 -90 7190
rect -30 6950 150 7190
rect 210 6950 390 7190
rect 450 6950 630 7190
rect 690 6950 1350 7190
rect 1410 6950 1430 7190
rect -360 6930 1430 6950
rect 2290 7190 4070 7210
rect 2290 6950 2310 7190
rect 2370 6950 3030 7190
rect 3090 6950 3270 7190
rect 3330 6950 3510 7190
rect 3570 6950 3750 7190
rect 3810 6950 3990 7190
rect 4050 6950 4070 7190
rect 2290 6930 4070 6950
rect 120 6220 240 6930
rect 1820 6640 1900 6660
rect 1820 6600 1840 6640
rect 1880 6600 1900 6640
rect 720 6360 810 6380
rect 720 6320 740 6360
rect 780 6320 810 6360
rect 720 6220 810 6320
rect 1440 6360 1530 6380
rect 1440 6320 1460 6360
rect 1500 6320 1530 6360
rect 1440 6220 1530 6320
rect -350 6200 -250 6220
rect -350 5960 -330 6200
rect -270 5960 -250 6200
rect -350 5940 -250 5960
rect -110 6200 470 6220
rect -110 5960 -90 6200
rect -30 5960 390 6200
rect 450 5960 470 6200
rect -110 5940 470 5960
rect 120 5930 470 5940
rect 710 6200 1570 6220
rect 710 5960 1350 6200
rect 1410 5960 1570 6200
rect 710 5940 1570 5960
rect 120 5380 240 5930
rect 710 5770 810 5940
rect 470 5740 810 5770
rect 470 5560 500 5740
rect 680 5560 810 5740
rect 470 5530 810 5560
rect 840 5460 1200 5510
rect 840 5380 930 5460
rect -350 5280 930 5380
rect 1110 5280 1200 5460
rect 1820 5430 1900 6600
rect 2050 6560 2150 6590
rect 2050 6520 2080 6560
rect 2120 6520 2150 6560
rect 2050 5750 2150 6520
rect 2190 6360 2280 6380
rect 2190 6320 2220 6360
rect 2260 6320 2280 6360
rect 2190 6220 2280 6320
rect 2900 6360 3000 6380
rect 2900 6320 2940 6360
rect 2980 6320 3000 6360
rect 2900 6220 3000 6320
rect 3480 6220 3600 6930
rect 5230 6430 5340 6450
rect 5230 6360 5250 6430
rect 5320 6360 5340 6430
rect 5230 6340 5340 6360
rect 2190 6200 3000 6220
rect 2190 5960 2310 6200
rect 2370 5960 3000 6200
rect 2190 5940 3000 5960
rect 3250 6200 3830 6220
rect 3250 5960 3270 6200
rect 3330 5960 3750 6200
rect 3810 5960 3830 6200
rect 3250 5940 3830 5960
rect 3970 6200 4120 6220
rect 3970 5960 3990 6200
rect 4050 5960 4120 6200
rect 3970 5940 4120 5960
rect 2050 5700 2070 5750
rect 2130 5700 2150 5750
rect 2050 5680 2150 5700
rect 2900 5770 3000 5940
rect 2900 5740 3270 5770
rect 2900 5560 3060 5740
rect 3240 5560 3270 5740
rect 2900 5530 3270 5560
rect 1820 5390 1840 5430
rect 1880 5390 1900 5430
rect 1820 5370 1900 5390
rect 2520 5460 2880 5510
rect 2520 5280 2610 5460
rect 2790 5410 2880 5460
rect 3480 5410 3600 5940
rect 2790 5320 4190 5410
rect 2790 5310 4070 5320
rect 2790 5280 3000 5310
rect -350 5130 -240 5280
rect 720 5240 1200 5280
rect 720 5200 760 5240
rect 800 5200 1200 5240
rect 720 5160 1200 5200
rect 1440 5240 1560 5280
rect 1440 5200 1480 5240
rect 1520 5200 1560 5240
rect 1440 5160 1560 5200
rect 2160 5240 2280 5280
rect 2160 5200 2200 5240
rect 2240 5200 2280 5240
rect 2160 5160 2280 5200
rect 2520 5270 3000 5280
rect 2520 5230 2920 5270
rect 2960 5230 3000 5270
rect 2520 5160 3000 5230
rect -350 4890 -330 5130
rect -270 4890 -240 5130
rect -350 4870 -240 4890
rect -110 5130 -10 5150
rect -110 4890 -90 5130
rect -30 4890 -10 5130
rect -110 4870 -10 4890
rect 370 5130 470 5150
rect 370 4890 390 5130
rect 450 4890 470 5130
rect 370 4870 470 4890
rect 720 5130 3000 5160
rect 720 4890 870 5130
rect 930 4890 2790 5130
rect 2850 4890 3000 5130
rect 720 4860 3000 4890
rect 3250 5130 3350 5150
rect 3250 4890 3270 5130
rect 3330 4890 3350 5130
rect 3250 4870 3350 4890
rect 3730 5130 3830 5150
rect 3730 4890 3750 5130
rect 3810 4890 3830 5130
rect 3730 4870 3830 4890
rect 3960 5130 4070 5310
rect 3960 4890 3990 5130
rect 4050 4890 4070 5130
rect 3960 4870 4070 4890
<< via1 >>
rect 3990 10000 4050 10010
rect 3990 9960 4000 10000
rect 4000 9960 4040 10000
rect 4040 9960 4050 10000
rect 3990 9950 4050 9960
rect 1240 9750 1300 9760
rect 1240 9710 1250 9750
rect 1250 9710 1290 9750
rect 1290 9710 1300 9750
rect 1240 9700 1300 9710
rect 2420 9750 2480 9760
rect 2420 9710 2430 9750
rect 2430 9710 2470 9750
rect 2470 9710 2480 9750
rect 2420 9700 2480 9710
rect -330 9380 -270 9620
rect -90 9380 -30 9620
rect 150 9380 210 9620
rect 390 9380 450 9620
rect 630 9380 690 9620
rect 1830 9380 1890 9620
rect 3030 9380 3090 9620
rect 3270 9380 3330 9620
rect 3510 9380 3570 9620
rect 3750 9380 3810 9620
rect 3990 9380 4050 9620
rect 730 9130 790 9190
rect -330 7830 -270 8070
rect -90 7830 -30 8070
rect 150 7830 210 8070
rect 390 7830 450 8070
rect 630 7830 690 8070
rect 1350 7830 1410 8070
rect 750 7600 810 7670
rect 2950 9130 3010 9190
rect 2310 7830 2370 8070
rect 3030 7830 3090 8070
rect 3270 7830 3330 8070
rect 3510 7830 3570 8070
rect 3750 7830 3810 8070
rect 3990 7830 4050 8070
rect 2910 7580 2970 7650
rect -330 5960 -270 6200
rect 500 5560 680 5740
rect 5250 6420 5320 6430
rect 5250 6370 5260 6420
rect 5260 6370 5310 6420
rect 5310 6370 5320 6420
rect 5250 6360 5320 6370
rect 3990 5960 4050 6200
rect 3060 5560 3240 5740
rect -90 4890 -30 5130
rect 390 4890 450 5130
rect 3270 4890 3330 5130
rect 3750 4890 3810 5130
<< metal2 >>
rect 3980 10010 4060 10020
rect 3980 9950 3990 10010
rect 4050 9950 4060 10010
rect 3980 9940 4060 9950
rect 1210 9760 1310 9780
rect 1210 9700 1240 9760
rect 1300 9700 1310 9760
rect 1210 9640 1310 9700
rect 2410 9760 2510 9780
rect 2410 9700 2420 9760
rect 2480 9700 2510 9760
rect 2410 9670 2510 9700
rect 2400 9640 2520 9670
rect -360 9620 4080 9640
rect -360 9380 -330 9620
rect -270 9380 -90 9620
rect -30 9380 150 9620
rect 210 9380 390 9620
rect 450 9380 630 9620
rect 690 9380 1830 9620
rect 1890 9380 3030 9620
rect 3090 9380 3270 9620
rect 3330 9380 3510 9620
rect 3570 9380 3750 9620
rect 3810 9380 3990 9620
rect 4050 9380 4080 9620
rect -360 9360 4080 9380
rect 1210 9210 1310 9360
rect 1810 9210 1910 9360
rect 2400 9210 2520 9360
rect 610 9190 3110 9210
rect 610 9130 730 9190
rect 790 9130 2950 9190
rect 3010 9130 3110 9190
rect 610 9110 3110 9130
rect 610 9100 820 9110
rect 2920 9100 3110 9110
rect 610 8090 710 9100
rect 3010 8090 3110 9100
rect -350 8070 1430 8090
rect -350 7830 -330 8070
rect -270 7830 -90 8070
rect -30 7830 150 8070
rect 210 7830 390 8070
rect 450 7830 630 8070
rect 690 7830 1350 8070
rect 1410 7830 1430 8070
rect -350 7810 1430 7830
rect 2290 8070 4070 8090
rect 2290 7830 2310 8070
rect 2370 7830 3030 8070
rect 3090 7830 3270 8070
rect 3330 7830 3510 8070
rect 3570 7830 3750 8070
rect 3810 7830 3990 8070
rect 4050 7830 4070 8070
rect 2290 7810 4070 7830
rect -350 6200 -250 7810
rect 710 7670 850 7810
rect 710 7600 750 7670
rect 810 7600 850 7670
rect 710 7520 850 7600
rect 2890 7650 2990 7810
rect 2890 7580 2910 7650
rect 2970 7580 2990 7650
rect 2890 7500 2990 7580
rect -350 5960 -330 6200
rect -270 5960 -250 6200
rect -350 5630 -250 5960
rect 3970 6200 4070 7810
rect 5230 6430 5340 6450
rect 5230 6360 5250 6430
rect 5320 6360 5340 6430
rect 5230 6340 5340 6360
rect 3970 5960 3990 6200
rect 4050 5960 4070 6200
rect 360 5740 710 5770
rect 360 5630 500 5740
rect -350 5560 500 5630
rect 680 5560 710 5740
rect -350 5530 710 5560
rect 3030 5740 3350 5770
rect 3030 5560 3060 5740
rect 3240 5630 3350 5740
rect 3970 5630 4070 5960
rect 3240 5560 4070 5630
rect 3030 5530 4070 5560
rect 360 5150 480 5530
rect -120 5130 480 5150
rect -120 4890 -90 5130
rect -30 4890 390 5130
rect 450 4890 480 5130
rect -120 4870 480 4890
rect 3250 5150 3350 5530
rect 3250 5130 3840 5150
rect 3250 4890 3270 5130
rect 3330 4890 3750 5130
rect 3810 4890 3840 5130
rect 3250 4870 3840 4890
<< via2 >>
rect 3990 9950 4050 10010
rect 5250 6360 5320 6430
<< metal3 >>
rect 3970 10020 4070 10030
rect 3970 9940 3980 10020
rect 4060 9940 4070 10020
rect 3970 9930 4070 9940
rect 5230 6430 5340 6490
rect 5230 6360 5250 6430
rect 5320 6360 5340 6430
rect 5230 6340 5340 6360
<< via3 >>
rect 3980 10010 4060 10020
rect 3980 9950 3990 10010
rect 3990 9950 4050 10010
rect 4050 9950 4060 10010
rect 3980 9940 4060 9950
<< metal4 >>
rect 3970 10020 4620 10030
rect 3970 9940 3980 10020
rect 4060 9940 4620 10020
rect 3970 9930 4620 9940
use sky130_fd_pr__cap_mim_m3_1_BW93LE  sky130_fd_pr__cap_mim_m3_1_BW93LE_0
timestamp 1620682856
transform 1 0 6780 0 1 8780
box -2350 -2300 2349 2300
use inverter_large  inverter_large_0
timestamp 1620670333
transform 1 0 4350 0 1 5520
box -240 -200 820 820
<< labels >>
rlabel poly -500 8400 -500 8400 7 VP
rlabel poly -500 9850 -500 9850 7 VN
rlabel locali 5420 5800 5420 5800 3 Vout
<< end >>
