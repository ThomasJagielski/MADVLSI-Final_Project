module decimation_filter (data_en,
    mclk1,
    mdata1,
    reset,
    VPWR,
    VGND,
    DATA,
    dec_rate);
 output data_en;
 input mclk1;
 input mdata1;
 input reset;
 input VPWR;
 input VGND;
 output [15:0] DATA;
 input [15:0] dec_rate;

 sky130_fd_sc_hd__or2_1 _2386_ (.A(_1891_),
    .B(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__or2_1 _2387_ (.A(_1826_),
    .B(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__a21oi_2 _2388_ (.A1(\acc3[23] ),
    .A2(\acc2[23] ),
    .B1(_1818_),
    .Y(_1896_));
 sky130_fd_sc_hd__inv_2 _2389_ (.A(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__o22a_1 _2390_ (.A1(\acc3[22] ),
    .A2(\acc2[22] ),
    .B1(_1540_),
    .B2(_0517_),
    .X(_1898_));
 sky130_fd_sc_hd__or4b_4 _2391_ (.A(_1895_),
    .B(_1897_),
    .C(_1823_),
    .D_N(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__o22a_2 _2392_ (.A1(_1818_),
    .A2(_1835_),
    .B1(_1889_),
    .B2(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__a22o_1 _2393_ (.A1(\acc3[28] ),
    .A2(\acc2[28] ),
    .B1(_1667_),
    .B2(_2350_),
    .X(_1901_));
 sky130_fd_sc_hd__o21ai_1 _2394_ (.A1(_1667_),
    .A2(_2350_),
    .B1(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hd__a22o_1 _2395_ (.A1(_1527_),
    .A2(_0504_),
    .B1(\acc3[24] ),
    .B2(\acc2[24] ),
    .X(_1903_));
 sky130_fd_sc_hd__o21ai_2 _2396_ (.A1(_1527_),
    .A2(_0504_),
    .B1(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__a211o_1 _2397_ (.A1(_1670_),
    .A2(_2366_),
    .B1(_1673_),
    .C1(_0499_),
    .X(_1905_));
 sky130_fd_sc_hd__o221a_1 _2398_ (.A1(_1670_),
    .A2(_2366_),
    .B1(_1811_),
    .B2(_1904_),
    .C1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__o32a_1 _2399_ (.A1(_1676_),
    .A2(_2358_),
    .A3(_1805_),
    .B1(_1677_),
    .B2(_0665_),
    .X(_1907_));
 sky130_fd_sc_hd__o221a_1 _2400_ (.A1(_1807_),
    .A2(_1902_),
    .B1(_1808_),
    .B2(_1906_),
    .C1(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__o31a_1 _2401_ (.A1(_1808_),
    .A2(_1817_),
    .A3(_1900_),
    .B1(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__o32a_1 _2402_ (.A1(_1681_),
    .A2(_2343_),
    .A3(_1794_),
    .B1(_1682_),
    .B2(_0670_),
    .X(_1910_));
 sky130_fd_sc_hd__o31a_1 _2403_ (.A1(_1796_),
    .A2(_1798_),
    .A3(_1909_),
    .B1(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__o32a_1 _2404_ (.A1(_1685_),
    .A2(_2335_),
    .A3(_1789_),
    .B1(_1686_),
    .B2(_0674_),
    .X(_1912_));
 sky130_fd_sc_hd__o31a_1 _2405_ (.A1(_1791_),
    .A2(_1793_),
    .A3(_1911_),
    .B1(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__inv_2 _2406_ (.A(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__inv_2 _2407_ (.A(_1788_),
    .Y(_1915_));
 sky130_fd_sc_hd__o221a_1 _2408_ (.A1(_1788_),
    .A2(_1914_),
    .B1(_1915_),
    .B2(_1913_),
    .C1(_1763_),
    .X(_0183_));
 sky130_fd_sc_hd__buf_1 _2409_ (.A(_0846_),
    .X(_1916_));
 sky130_fd_sc_hd__buf_1 _2410_ (.A(_1916_),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _2411_ (.A(_1911_),
    .B(_1793_),
    .X(_1917_));
 sky130_fd_sc_hd__o21ai_1 _2412_ (.A1(_1685_),
    .A2(_2335_),
    .B1(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__inv_2 _2413_ (.A(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__o221a_1 _2414_ (.A1(_1791_),
    .A2(_1919_),
    .B1(_1790_),
    .B2(_1918_),
    .C1(_1763_),
    .X(_0182_));
 sky130_fd_sc_hd__buf_1 _2415_ (.A(_1916_),
    .X(_0070_));
 sky130_fd_sc_hd__inv_2 _2416_ (.A(_1911_),
    .Y(_1920_));
 sky130_fd_sc_hd__clkbuf_2 _2417_ (.A(_0687_),
    .X(_1921_));
 sky130_fd_sc_hd__o211a_1 _2418_ (.A1(_1920_),
    .A2(_1792_),
    .B1(_1921_),
    .C1(_1917_),
    .X(_0181_));
 sky130_fd_sc_hd__buf_1 _2419_ (.A(_1916_),
    .X(_0069_));
 sky130_fd_sc_hd__or2_1 _2420_ (.A(_1909_),
    .B(_1798_),
    .X(_1922_));
 sky130_fd_sc_hd__o21ai_1 _2421_ (.A1(_1681_),
    .A2(_2343_),
    .B1(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__inv_2 _2422_ (.A(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__buf_2 _2423_ (.A(_1708_),
    .X(_1925_));
 sky130_fd_sc_hd__o221a_1 _2424_ (.A1(_1796_),
    .A2(_1924_),
    .B1(_1795_),
    .B2(_1923_),
    .C1(_1925_),
    .X(_0180_));
 sky130_fd_sc_hd__buf_1 _2425_ (.A(_1916_),
    .X(_0068_));
 sky130_fd_sc_hd__inv_2 _2426_ (.A(_1909_),
    .Y(_1926_));
 sky130_fd_sc_hd__o211a_1 _2427_ (.A1(_1926_),
    .A2(_1797_),
    .B1(_1921_),
    .C1(_1922_),
    .X(_0179_));
 sky130_fd_sc_hd__buf_1 _2428_ (.A(_1916_),
    .X(_0067_));
 sky130_fd_sc_hd__o21ai_1 _2429_ (.A1(_1900_),
    .A2(_1817_),
    .B1(_1906_),
    .Y(_1927_));
 sky130_fd_sc_hd__inv_2 _2430_ (.A(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__o21ai_1 _2431_ (.A1(_1803_),
    .A2(_1928_),
    .B1(_1902_),
    .Y(_1929_));
 sky130_fd_sc_hd__nand2_1 _2432_ (.A(_1804_),
    .B(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__o21ai_1 _2433_ (.A1(_1676_),
    .A2(_2358_),
    .B1(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _2434_ (.A(_1806_),
    .B(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__o211a_1 _2435_ (.A1(_1806_),
    .A2(_1931_),
    .B1(_1921_),
    .C1(_1932_),
    .X(_0178_));
 sky130_fd_sc_hd__buf_1 _2436_ (.A(_0846_),
    .X(_1933_));
 sky130_fd_sc_hd__buf_1 _2437_ (.A(_1933_),
    .X(_0066_));
 sky130_fd_sc_hd__o211a_1 _2438_ (.A1(_1804_),
    .A2(_1929_),
    .B1(_1921_),
    .C1(_1930_),
    .X(_0177_));
 sky130_fd_sc_hd__buf_1 _2439_ (.A(_1933_),
    .X(_0065_));
 sky130_fd_sc_hd__or2_1 _2440_ (.A(_1800_),
    .B(_1928_),
    .X(_1934_));
 sky130_fd_sc_hd__o21ai_1 _2441_ (.A1(_1506_),
    .A2(_2347_),
    .B1(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__inv_2 _2442_ (.A(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__o221a_1 _2443_ (.A1(_1802_),
    .A2(_1936_),
    .B1(_1801_),
    .B2(_1935_),
    .C1(_1925_),
    .X(_0176_));
 sky130_fd_sc_hd__buf_1 _2444_ (.A(_1933_),
    .X(_0064_));
 sky130_fd_sc_hd__o211a_1 _2445_ (.A1(_1799_),
    .A2(_1927_),
    .B1(_1921_),
    .C1(_1934_),
    .X(_0175_));
 sky130_fd_sc_hd__buf_1 _2446_ (.A(_1933_),
    .X(_0063_));
 sky130_fd_sc_hd__o21ai_1 _2447_ (.A1(_1900_),
    .A2(_1816_),
    .B1(_1904_),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _2448_ (.A(_1810_),
    .B(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__o21ai_1 _2449_ (.A1(_1673_),
    .A2(_0499_),
    .B1(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__buf_2 _2450_ (.A(_0687_),
    .X(_1940_));
 sky130_fd_sc_hd__nand2_1 _2451_ (.A(_1809_),
    .B(_1939_),
    .Y(_1941_));
 sky130_fd_sc_hd__o211a_1 _2452_ (.A1(_1809_),
    .A2(_1939_),
    .B1(_1940_),
    .C1(_1941_),
    .X(_0174_));
 sky130_fd_sc_hd__buf_1 _2453_ (.A(_1933_),
    .X(_0062_));
 sky130_fd_sc_hd__o211a_1 _2454_ (.A1(_1810_),
    .A2(_1937_),
    .B1(_1940_),
    .C1(_1938_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_1 _2455_ (.A(_0846_),
    .X(_1942_));
 sky130_fd_sc_hd__buf_1 _2456_ (.A(_1942_),
    .X(_0061_));
 sky130_fd_sc_hd__or2_1 _2457_ (.A(_1900_),
    .B(_1815_),
    .X(_1943_));
 sky130_fd_sc_hd__o21ai_1 _2458_ (.A1(_1532_),
    .A2(_0508_),
    .B1(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__inv_2 _2459_ (.A(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__o221a_1 _2460_ (.A1(_1813_),
    .A2(_1945_),
    .B1(_1812_),
    .B2(_1944_),
    .C1(_1925_),
    .X(_0172_));
 sky130_fd_sc_hd__buf_1 _2461_ (.A(_1942_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _2462_ (.A(_1900_),
    .Y(_1946_));
 sky130_fd_sc_hd__o211a_1 _2463_ (.A1(_1946_),
    .A2(_1814_),
    .B1(_1940_),
    .C1(_1943_),
    .X(_0171_));
 sky130_fd_sc_hd__buf_1 _2464_ (.A(_1942_),
    .X(_0059_));
 sky130_fd_sc_hd__o21ai_1 _2465_ (.A1(_1889_),
    .A2(_1895_),
    .B1(_1830_),
    .Y(_1947_));
 sky130_fd_sc_hd__inv_2 _2466_ (.A(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__o21ai_1 _2467_ (.A1(_1823_),
    .A2(_1948_),
    .B1(_1833_),
    .Y(_1949_));
 sky130_fd_sc_hd__nand2_1 _2468_ (.A(_1898_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__o21ai_1 _2469_ (.A1(_1541_),
    .A2(_0518_),
    .B1(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hd__inv_2 _2470_ (.A(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__o221a_1 _2471_ (.A1(_1897_),
    .A2(_1952_),
    .B1(_1896_),
    .B2(_1951_),
    .C1(_1925_),
    .X(_0170_));
 sky130_fd_sc_hd__buf_1 _2472_ (.A(_1942_),
    .X(_0058_));
 sky130_fd_sc_hd__o211a_1 _2473_ (.A1(_1898_),
    .A2(_1949_),
    .B1(_1940_),
    .C1(_1950_),
    .X(_0169_));
 sky130_fd_sc_hd__buf_1 _2474_ (.A(_1942_),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _2475_ (.A(_1822_),
    .B(_1948_),
    .X(_1953_));
 sky130_fd_sc_hd__o21ai_1 _2476_ (.A1(_1548_),
    .A2(_0525_),
    .B1(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__inv_2 _2477_ (.A(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__o221a_1 _2478_ (.A1(_1820_),
    .A2(_1955_),
    .B1(_1819_),
    .B2(_1954_),
    .C1(_1925_),
    .X(_0168_));
 sky130_fd_sc_hd__buf_1 _2479_ (.A(_0846_),
    .X(_1956_));
 sky130_fd_sc_hd__buf_1 _2480_ (.A(_1956_),
    .X(_0056_));
 sky130_fd_sc_hd__o211a_1 _2481_ (.A1(_1821_),
    .A2(_1947_),
    .B1(_1940_),
    .C1(_1953_),
    .X(_0167_));
 sky130_fd_sc_hd__buf_1 _2482_ (.A(_1956_),
    .X(_0055_));
 sky130_fd_sc_hd__o21ai_1 _2483_ (.A1(_1889_),
    .A2(_1894_),
    .B1(_1828_),
    .Y(_1957_));
 sky130_fd_sc_hd__nand2_1 _2484_ (.A(_1825_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__o21ai_1 _2485_ (.A1(_1563_),
    .A2(_0535_),
    .B1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__clkbuf_2 _2486_ (.A(_0687_),
    .X(_1960_));
 sky130_fd_sc_hd__nand2_1 _2487_ (.A(_1824_),
    .B(_1959_),
    .Y(_1961_));
 sky130_fd_sc_hd__o211a_1 _2488_ (.A1(_1824_),
    .A2(_1959_),
    .B1(_1960_),
    .C1(_1961_),
    .X(_0166_));
 sky130_fd_sc_hd__buf_1 _2489_ (.A(_1956_),
    .X(_0054_));
 sky130_fd_sc_hd__o211a_1 _2490_ (.A1(_1825_),
    .A2(_1957_),
    .B1(_1960_),
    .C1(_1958_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_1 _2491_ (.A(_1956_),
    .X(_0053_));
 sky130_fd_sc_hd__or2_1 _2492_ (.A(_1889_),
    .B(_1893_),
    .X(_1962_));
 sky130_fd_sc_hd__o21ai_1 _2493_ (.A1(_1657_),
    .A2(_0648_),
    .B1(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__inv_2 _2494_ (.A(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__buf_2 _2495_ (.A(_1708_),
    .X(_1965_));
 sky130_fd_sc_hd__o221a_1 _2496_ (.A1(_1891_),
    .A2(_1964_),
    .B1(_1890_),
    .B2(_1963_),
    .C1(_1965_),
    .X(_0164_));
 sky130_fd_sc_hd__buf_1 _2497_ (.A(_1956_),
    .X(_0052_));
 sky130_fd_sc_hd__inv_2 _2498_ (.A(_1889_),
    .Y(_1966_));
 sky130_fd_sc_hd__o211a_1 _2499_ (.A1(_1966_),
    .A2(_1892_),
    .B1(_1960_),
    .C1(_1962_),
    .X(_0163_));
 sky130_fd_sc_hd__buf_1 _2500_ (.A(_0734_),
    .X(_1967_));
 sky130_fd_sc_hd__buf_1 _2501_ (.A(_1967_),
    .X(_0051_));
 sky130_fd_sc_hd__o21ai_1 _2502_ (.A1(_1880_),
    .A2(_1854_),
    .B1(_1886_),
    .Y(_1968_));
 sky130_fd_sc_hd__inv_2 _2503_ (.A(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__o21ai_1 _2504_ (.A1(_1844_),
    .A2(_1969_),
    .B1(_1882_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _2505_ (.A(_1838_),
    .B(_1970_),
    .Y(_1971_));
 sky130_fd_sc_hd__o21ai_1 _2506_ (.A1(_1649_),
    .A2(_0552_),
    .B1(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__nand2_1 _2507_ (.A(_1837_),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__o211a_1 _2508_ (.A1(_1837_),
    .A2(_1972_),
    .B1(_1960_),
    .C1(_1973_),
    .X(_0162_));
 sky130_fd_sc_hd__buf_1 _2509_ (.A(_1967_),
    .X(_0050_));
 sky130_fd_sc_hd__o211a_1 _2510_ (.A1(_1838_),
    .A2(_1970_),
    .B1(_1960_),
    .C1(_1971_),
    .X(_0161_));
 sky130_fd_sc_hd__buf_1 _2511_ (.A(_1967_),
    .X(_0049_));
 sky130_fd_sc_hd__or2_1 _2512_ (.A(_1843_),
    .B(_1969_),
    .X(_1974_));
 sky130_fd_sc_hd__o21ai_1 _2513_ (.A1(_1584_),
    .A2(_0561_),
    .B1(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__inv_2 _2514_ (.A(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__o221a_1 _2515_ (.A1(_1841_),
    .A2(_1976_),
    .B1(_1840_),
    .B2(_1975_),
    .C1(_1965_),
    .X(_0160_));
 sky130_fd_sc_hd__buf_1 _2516_ (.A(_1967_),
    .X(_0048_));
 sky130_fd_sc_hd__clkbuf_2 _2517_ (.A(_0687_),
    .X(_1977_));
 sky130_fd_sc_hd__o211a_1 _2518_ (.A1(_1842_),
    .A2(_1968_),
    .B1(_1977_),
    .C1(_1974_),
    .X(_0159_));
 sky130_fd_sc_hd__buf_1 _2519_ (.A(_1967_),
    .X(_0047_));
 sky130_fd_sc_hd__o21ai_1 _2520_ (.A1(_1880_),
    .A2(_1853_),
    .B1(_1884_),
    .Y(_1978_));
 sky130_fd_sc_hd__nand2_1 _2521_ (.A(_1847_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__o21ai_1 _2522_ (.A1(_1646_),
    .A2(_0572_),
    .B1(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _2523_ (.A(_1846_),
    .B(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__o211a_1 _2524_ (.A1(_1846_),
    .A2(_1980_),
    .B1(_1977_),
    .C1(_1981_),
    .X(_0158_));
 sky130_fd_sc_hd__buf_1 _2525_ (.A(_0734_),
    .X(_1982_));
 sky130_fd_sc_hd__buf_1 _2526_ (.A(_1982_),
    .X(_0046_));
 sky130_fd_sc_hd__o211a_1 _2527_ (.A1(_1847_),
    .A2(_1978_),
    .B1(_1977_),
    .C1(_1979_),
    .X(_0157_));
 sky130_fd_sc_hd__buf_1 _2528_ (.A(_1982_),
    .X(_0045_));
 sky130_fd_sc_hd__or2_1 _2529_ (.A(_1880_),
    .B(_1852_),
    .X(_1983_));
 sky130_fd_sc_hd__o21ai_1 _2530_ (.A1(_1599_),
    .A2(_0581_),
    .B1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__inv_2 _2531_ (.A(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hd__o221a_1 _2532_ (.A1(_1850_),
    .A2(_1985_),
    .B1(_1849_),
    .B2(_1984_),
    .C1(_1965_),
    .X(_0156_));
 sky130_fd_sc_hd__buf_1 _2533_ (.A(_1982_),
    .X(_0044_));
 sky130_fd_sc_hd__inv_2 _2534_ (.A(_1880_),
    .Y(_1986_));
 sky130_fd_sc_hd__o211a_1 _2535_ (.A1(_1986_),
    .A2(_1851_),
    .B1(_1977_),
    .C1(_1983_),
    .X(_0155_));
 sky130_fd_sc_hd__buf_1 _2536_ (.A(_1982_),
    .X(_0043_));
 sky130_fd_sc_hd__inv_2 _2537_ (.A(_1878_),
    .Y(_1987_));
 sky130_fd_sc_hd__a31o_1 _2538_ (.A1(_1865_),
    .A2(_1866_),
    .A3(_1987_),
    .B1(_1862_),
    .X(_1988_));
 sky130_fd_sc_hd__nand2_1 _2539_ (.A(_1858_),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__o21ai_1 _2540_ (.A1(_1616_),
    .A2(_0591_),
    .B1(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__inv_2 _2541_ (.A(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__o221a_1 _2542_ (.A1(_1857_),
    .A2(_1991_),
    .B1(_1856_),
    .B2(_1990_),
    .C1(_1965_),
    .X(_0154_));
 sky130_fd_sc_hd__buf_1 _2543_ (.A(_1982_),
    .X(_0042_));
 sky130_fd_sc_hd__o211a_1 _2544_ (.A1(_1858_),
    .A2(_1988_),
    .B1(_1977_),
    .C1(_1989_),
    .X(_0153_));
 sky130_fd_sc_hd__buf_1 _2545_ (.A(_0734_),
    .X(_1992_));
 sky130_fd_sc_hd__buf_1 _2546_ (.A(_1992_),
    .X(_0041_));
 sky130_fd_sc_hd__nand2_1 _2547_ (.A(_1987_),
    .B(_1866_),
    .Y(_1993_));
 sky130_fd_sc_hd__inv_2 _2548_ (.A(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__o21ai_1 _2549_ (.A1(_1861_),
    .A2(_1994_),
    .B1(_1865_),
    .Y(_1995_));
 sky130_fd_sc_hd__o311a_1 _2550_ (.A1(_1861_),
    .A2(_1994_),
    .A3(_1865_),
    .B1(_0688_),
    .C1(_1995_),
    .X(_0152_));
 sky130_fd_sc_hd__buf_1 _2551_ (.A(_1992_),
    .X(_0040_));
 sky130_fd_sc_hd__o211a_1 _2552_ (.A1(_1987_),
    .A2(_1866_),
    .B1(_0774_),
    .C1(_1993_),
    .X(_0151_));
 sky130_fd_sc_hd__buf_1 _2553_ (.A(_1992_),
    .X(_0039_));
 sky130_fd_sc_hd__or2_1 _2554_ (.A(_1876_),
    .B(_1872_),
    .X(_1996_));
 sky130_fd_sc_hd__o21ai_1 _2555_ (.A1(_1635_),
    .A2(_0613_),
    .B1(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__inv_2 _2556_ (.A(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__o221a_1 _2557_ (.A1(_1870_),
    .A2(_1998_),
    .B1(_1869_),
    .B2(_1997_),
    .C1(_1965_),
    .X(_0150_));
 sky130_fd_sc_hd__buf_1 _2558_ (.A(_1992_),
    .X(_0038_));
 sky130_fd_sc_hd__o211a_1 _2559_ (.A1(_1875_),
    .A2(_1871_),
    .B1(_0774_),
    .C1(_1996_),
    .X(_0149_));
 sky130_fd_sc_hd__buf_1 _2560_ (.A(_1992_),
    .X(_0037_));
 sky130_fd_sc_hd__o21a_1 _2561_ (.A1(_1778_),
    .A2(_0621_),
    .B1(_1873_),
    .X(_1999_));
 sky130_fd_sc_hd__and3b_1 _2562_ (.A_N(_1999_),
    .B(_1874_),
    .C(_0774_),
    .X(_0148_));
 sky130_fd_sc_hd__buf_1 _2563_ (.A(_2326_),
    .X(_0036_));
 sky130_fd_sc_hd__o221a_1 _2564_ (.A1(_1778_),
    .A2(_0621_),
    .B1(\acc3[0] ),
    .B2(\acc2[0] ),
    .C1(_1173_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_2 _2565_ (.A(\diff3[8] ),
    .X(_2000_));
 sky130_fd_sc_hd__or2_2 _2566_ (.A(\diff3[13] ),
    .B(\diff3[12] ),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_2 _2567_ (.A(\diff3[24] ),
    .X(_2002_));
 sky130_fd_sc_hd__or3b_1 _2568_ (.A(\diff3[19] ),
    .B(\diff3[18] ),
    .C_N(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__or4_4 _2569_ (.A(\diff3[21] ),
    .B(\diff3[23] ),
    .C(\diff3[22] ),
    .D(\diff3[20] ),
    .X(_2004_));
 sky130_fd_sc_hd__or4_4 _2570_ (.A(\diff3[14] ),
    .B(\diff3[15] ),
    .C(\diff3[17] ),
    .D(\diff3[16] ),
    .X(_2005_));
 sky130_fd_sc_hd__or4_4 _2571_ (.A(\diff3[9] ),
    .B(\diff3[8] ),
    .C(\diff3[11] ),
    .D(\diff3[10] ),
    .X(_2006_));
 sky130_fd_sc_hd__or2_1 _2572_ (.A(_2005_),
    .B(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__nor4_2 _2573_ (.A(_2001_),
    .B(_2003_),
    .C(_2004_),
    .D(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__buf_1 _2574_ (.A(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__or2_1 _2575_ (.A(_2000_),
    .B(_2009_),
    .X(_0032_));
 sky130_fd_sc_hd__or3_1 _2576_ (.A(_2266_),
    .B(net3),
    .C(_2257_),
    .X(_2010_));
 sky130_fd_sc_hd__or3_4 _2577_ (.A(net15),
    .B(net16),
    .C(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__nor3_4 _2578_ (.A(_2282_),
    .B(_2011_),
    .C(_0897_),
    .Y(_2012_));
 sky130_fd_sc_hd__buf_1 _2579_ (.A(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__or2_1 _2580_ (.A(net14),
    .B(_2011_),
    .X(_2014_));
 sky130_fd_sc_hd__or4_4 _2581_ (.A(_2312_),
    .B(_2292_),
    .C(_0895_),
    .D(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__inv_2 _2582_ (.A(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__clkbuf_2 _2583_ (.A(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__or3b_4 _2584_ (.A(_0896_),
    .B(_2014_),
    .C_N(_2292_),
    .X(_2018_));
 sky130_fd_sc_hd__inv_2 _2585_ (.A(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__clkbuf_2 _2586_ (.A(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__or4_4 _2587_ (.A(_0873_),
    .B(_2251_),
    .C(_0881_),
    .D(_2010_),
    .X(_2021_));
 sky130_fd_sc_hd__inv_2 _2588_ (.A(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__buf_1 _2589_ (.A(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__or4_4 _2590_ (.A(_2013_),
    .B(_2017_),
    .C(_2020_),
    .D(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__or4b_4 _2591_ (.A(_0883_),
    .B(net3),
    .C(_2257_),
    .D_N(_2266_),
    .X(_2025_));
 sky130_fd_sc_hd__or4_4 _2592_ (.A(net6),
    .B(net7),
    .C(_0886_),
    .D(net5),
    .X(_2026_));
 sky130_fd_sc_hd__or3_4 _2593_ (.A(_0873_),
    .B(_2258_),
    .C(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__or3_4 _2594_ (.A(_2265_),
    .B(_0892_),
    .C(_2257_),
    .X(_2028_));
 sky130_fd_sc_hd__and4b_4 _2595_ (.A_N(_2024_),
    .B(_2025_),
    .C(_2027_),
    .D(_2028_),
    .X(_0033_));
 sky130_fd_sc_hd__clkbuf_2 _2596_ (.A(\diff3[20] ),
    .X(_2029_));
 sky130_fd_sc_hd__or2_1 _2597_ (.A(\diff3[29] ),
    .B(\diff3[28] ),
    .X(_2030_));
 sky130_fd_sc_hd__or3_4 _2598_ (.A(\diff3[30] ),
    .B(\diff3[32] ),
    .C(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__or3b_2 _2599_ (.A(\diff3[35] ),
    .B(\diff3[34] ),
    .C_N(\diff3[36] ),
    .X(_2032_));
 sky130_fd_sc_hd__or3_4 _2600_ (.A(\diff3[31] ),
    .B(\diff3[33] ),
    .C(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__clkbuf_2 _2601_ (.A(\diff3[27] ),
    .X(_2034_));
 sky130_fd_sc_hd__or2_2 _2602_ (.A(\diff3[25] ),
    .B(\diff3[26] ),
    .X(_2035_));
 sky130_fd_sc_hd__or4_4 _2603_ (.A(\diff3[24] ),
    .B(_2034_),
    .C(_2035_),
    .D(_2004_),
    .X(_2036_));
 sky130_fd_sc_hd__nor3_4 _2604_ (.A(_2031_),
    .B(_2033_),
    .C(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__clkbuf_2 _2605_ (.A(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__nor2_1 _2606_ (.A(_2029_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__clkbuf_2 _2607_ (.A(\diff3[17] ),
    .X(_2040_));
 sky130_fd_sc_hd__or4_4 _2608_ (.A(\diff3[19] ),
    .B(\diff3[18] ),
    .C(\diff3[17] ),
    .D(\diff3[20] ),
    .X(_2041_));
 sky130_fd_sc_hd__or4_4 _2609_ (.A(\diff3[21] ),
    .B(\diff3[23] ),
    .C(\diff3[22] ),
    .D(\diff3[24] ),
    .X(_2042_));
 sky130_fd_sc_hd__or4b_4 _2610_ (.A(_2034_),
    .B(\diff3[31] ),
    .C(_2042_),
    .D_N(\diff3[33] ),
    .X(_2043_));
 sky130_fd_sc_hd__nor4_2 _2611_ (.A(_2031_),
    .B(_2035_),
    .C(_2041_),
    .D(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__clkbuf_2 _2612_ (.A(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__nor2_1 _2613_ (.A(_2040_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__clkbuf_2 _2614_ (.A(\diff3[14] ),
    .X(_2047_));
 sky130_fd_sc_hd__or4b_4 _2615_ (.A(\diff3[19] ),
    .B(\diff3[18] ),
    .C(_2030_),
    .D_N(\diff3[30] ),
    .X(_2048_));
 sky130_fd_sc_hd__nor3_4 _2616_ (.A(_2005_),
    .B(_2048_),
    .C(_2036_),
    .Y(_2049_));
 sky130_fd_sc_hd__nor2_1 _2617_ (.A(_2047_),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__clkbuf_2 _2618_ (.A(\diff3[11] ),
    .X(_2051_));
 sky130_fd_sc_hd__or3_1 _2619_ (.A(\diff3[11] ),
    .B(\diff3[15] ),
    .C(\diff3[16] ),
    .X(_2052_));
 sky130_fd_sc_hd__or4_4 _2620_ (.A(\diff3[14] ),
    .B(_2001_),
    .C(_2052_),
    .D(_2041_),
    .X(_2053_));
 sky130_fd_sc_hd__or4b_4 _2621_ (.A(_2053_),
    .B(_2035_),
    .C(_2042_),
    .D_N(\diff3[27] ),
    .X(_2054_));
 sky130_fd_sc_hd__inv_2 _2622_ (.A(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2623_ (.A(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__nor2_1 _2624_ (.A(_2051_),
    .B(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__or4_4 _2625_ (.A(\diff3[5] ),
    .B(\diff3[2] ),
    .C(\diff3[3] ),
    .D(\diff3[4] ),
    .X(_2058_));
 sky130_fd_sc_hd__or3_1 _2626_ (.A(\diff3[6] ),
    .B(\diff3[7] ),
    .C(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__or4b_4 _2627_ (.A(_2059_),
    .B(_2001_),
    .C(_2007_),
    .D_N(\diff3[18] ),
    .X(_2060_));
 sky130_fd_sc_hd__inv_2 _2628_ (.A(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__clkbuf_2 _2629_ (.A(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__nor2_1 _2630_ (.A(\diff3[2] ),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__or4b_4 _2631_ (.A(_2006_),
    .B(\diff3[1] ),
    .C(\diff3[0] ),
    .D_N(\diff3[15] ),
    .X(_2064_));
 sky130_fd_sc_hd__or4_4 _2632_ (.A(\diff3[14] ),
    .B(_2001_),
    .C(_2064_),
    .D(_2059_),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_2 _2633_ (.A(\diff3[10] ),
    .X(_2066_));
 sky130_fd_sc_hd__or2b_1 _2634_ (.A(_2066_),
    .B_N(\diff3[21] ),
    .X(_2067_));
 sky130_fd_sc_hd__clkbuf_2 _2635_ (.A(\diff3[9] ),
    .X(_2068_));
 sky130_fd_sc_hd__or4_4 _2636_ (.A(_2068_),
    .B(_2000_),
    .C(\diff3[6] ),
    .D(\diff3[7] ),
    .X(_2069_));
 sky130_fd_sc_hd__nor4_2 _2637_ (.A(\diff3[5] ),
    .B(_2067_),
    .C(_2069_),
    .D(_2053_),
    .Y(_2070_));
 sky130_fd_sc_hd__clkbuf_2 _2638_ (.A(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__o21ai_1 _2639_ (.A1(\diff3[5] ),
    .A2(_2071_),
    .B1(_2013_),
    .Y(_2072_));
 sky130_fd_sc_hd__o221a_1 _2640_ (.A1(_2018_),
    .A2(_2063_),
    .B1(_2015_),
    .B2(_2065_),
    .C1(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__o221a_1 _2641_ (.A1(_2025_),
    .A2(_2050_),
    .B1(_2021_),
    .B2(_2057_),
    .C1(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__o221ai_1 _2642_ (.A1(_2027_),
    .A2(_2039_),
    .B1(_2028_),
    .B2(_2046_),
    .C1(_2074_),
    .Y(_0034_));
 sky130_fd_sc_hd__or2_1 _2643_ (.A(_2068_),
    .B(_2009_),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_2 _2644_ (.A(\diff3[15] ),
    .X(_2075_));
 sky130_fd_sc_hd__buf_1 _2645_ (.A(_2049_),
    .X(_2076_));
 sky130_fd_sc_hd__inv_2 _2646_ (.A(_2025_),
    .Y(_2077_));
 sky130_fd_sc_hd__buf_1 _2647_ (.A(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__o21a_1 _2648_ (.A1(_2075_),
    .A2(_2076_),
    .B1(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__o21a_1 _2649_ (.A1(\diff3[6] ),
    .A2(_2071_),
    .B1(_2013_),
    .X(_2080_));
 sky130_fd_sc_hd__inv_2 _2650_ (.A(_2065_),
    .Y(_2081_));
 sky130_fd_sc_hd__clkbuf_2 _2651_ (.A(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__o21a_1 _2652_ (.A1(\diff3[0] ),
    .A2(_2082_),
    .B1(_2017_),
    .X(_2083_));
 sky130_fd_sc_hd__o21a_1 _2653_ (.A1(\diff3[3] ),
    .A2(_2062_),
    .B1(_2020_),
    .X(_2084_));
 sky130_fd_sc_hd__clkbuf_2 _2654_ (.A(\diff3[12] ),
    .X(_2085_));
 sky130_fd_sc_hd__o21a_1 _2655_ (.A1(_2085_),
    .A2(_2056_),
    .B1(_2023_),
    .X(_2086_));
 sky130_fd_sc_hd__or4_4 _2656_ (.A(_2080_),
    .B(_2083_),
    .C(_2084_),
    .D(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__clkbuf_2 _2657_ (.A(\diff3[21] ),
    .X(_2088_));
 sky130_fd_sc_hd__inv_2 _2658_ (.A(_2027_),
    .Y(_2089_));
 sky130_fd_sc_hd__buf_1 _2659_ (.A(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__o21a_1 _2660_ (.A1(_2088_),
    .A2(_2038_),
    .B1(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__clkbuf_2 _2661_ (.A(\diff3[18] ),
    .X(_2092_));
 sky130_fd_sc_hd__inv_2 _2662_ (.A(_2028_),
    .Y(_2093_));
 sky130_fd_sc_hd__buf_1 _2663_ (.A(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__o21a_1 _2664_ (.A1(_2092_),
    .A2(_2045_),
    .B1(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__or4_1 _2665_ (.A(_2079_),
    .B(_2087_),
    .C(_2091_),
    .D(_2095_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _2666_ (.A(_2066_),
    .B(_2009_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_2 _2667_ (.A(\diff3[16] ),
    .X(_2096_));
 sky130_fd_sc_hd__o21a_1 _2668_ (.A1(_2096_),
    .A2(_2076_),
    .B1(_2078_),
    .X(_2097_));
 sky130_fd_sc_hd__o21a_1 _2669_ (.A1(\diff3[7] ),
    .A2(_2071_),
    .B1(_2013_),
    .X(_2098_));
 sky130_fd_sc_hd__o21a_1 _2670_ (.A1(\diff3[1] ),
    .A2(_2082_),
    .B1(_2017_),
    .X(_2099_));
 sky130_fd_sc_hd__o21a_1 _2671_ (.A1(\diff3[4] ),
    .A2(_2062_),
    .B1(_2020_),
    .X(_2100_));
 sky130_fd_sc_hd__clkbuf_2 _2672_ (.A(\diff3[13] ),
    .X(_2101_));
 sky130_fd_sc_hd__o21a_1 _2673_ (.A1(_2101_),
    .A2(_2056_),
    .B1(_2023_),
    .X(_2102_));
 sky130_fd_sc_hd__or4_4 _2674_ (.A(_2098_),
    .B(_2099_),
    .C(_2100_),
    .D(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__clkbuf_2 _2675_ (.A(\diff3[22] ),
    .X(_2104_));
 sky130_fd_sc_hd__o21a_1 _2676_ (.A1(_2104_),
    .A2(_2038_),
    .B1(_2090_),
    .X(_2105_));
 sky130_fd_sc_hd__clkbuf_2 _2677_ (.A(\diff3[19] ),
    .X(_2106_));
 sky130_fd_sc_hd__o21a_1 _2678_ (.A1(_2106_),
    .A2(_2045_),
    .B1(_2094_),
    .X(_2107_));
 sky130_fd_sc_hd__or4_1 _2679_ (.A(_2097_),
    .B(_2103_),
    .C(_2105_),
    .D(_2107_),
    .X(_0003_));
 sky130_fd_sc_hd__or2_1 _2680_ (.A(_2051_),
    .B(_2009_),
    .X(_0004_));
 sky130_fd_sc_hd__o21a_1 _2681_ (.A1(_2040_),
    .A2(_2076_),
    .B1(_2078_),
    .X(_2108_));
 sky130_fd_sc_hd__o21a_1 _2682_ (.A1(_2000_),
    .A2(_2071_),
    .B1(_2013_),
    .X(_2109_));
 sky130_fd_sc_hd__o21a_1 _2683_ (.A1(\diff3[2] ),
    .A2(_2082_),
    .B1(_2017_),
    .X(_2110_));
 sky130_fd_sc_hd__o21a_1 _2684_ (.A1(\diff3[5] ),
    .A2(_2062_),
    .B1(_2020_),
    .X(_2111_));
 sky130_fd_sc_hd__o21a_1 _2685_ (.A1(_2047_),
    .A2(_2056_),
    .B1(_2023_),
    .X(_2112_));
 sky130_fd_sc_hd__or4_4 _2686_ (.A(_2109_),
    .B(_2110_),
    .C(_2111_),
    .D(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__clkbuf_2 _2687_ (.A(\diff3[23] ),
    .X(_2114_));
 sky130_fd_sc_hd__o21a_1 _2688_ (.A1(_2114_),
    .A2(_2038_),
    .B1(_2090_),
    .X(_2115_));
 sky130_fd_sc_hd__o21a_1 _2689_ (.A1(_2029_),
    .A2(_2045_),
    .B1(_2094_),
    .X(_2116_));
 sky130_fd_sc_hd__or4_1 _2690_ (.A(_2108_),
    .B(_2113_),
    .C(_2115_),
    .D(_2116_),
    .X(_0005_));
 sky130_fd_sc_hd__or2_1 _2691_ (.A(_2085_),
    .B(_2009_),
    .X(_0006_));
 sky130_fd_sc_hd__o21a_1 _2692_ (.A1(_2092_),
    .A2(_2076_),
    .B1(_2078_),
    .X(_2117_));
 sky130_fd_sc_hd__buf_1 _2693_ (.A(_2012_),
    .X(_2118_));
 sky130_fd_sc_hd__o21a_1 _2694_ (.A1(_2068_),
    .A2(_2071_),
    .B1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__o21a_1 _2695_ (.A1(\diff3[3] ),
    .A2(_2082_),
    .B1(_2017_),
    .X(_2120_));
 sky130_fd_sc_hd__o21a_1 _2696_ (.A1(\diff3[6] ),
    .A2(_2062_),
    .B1(_2020_),
    .X(_2121_));
 sky130_fd_sc_hd__o21a_1 _2697_ (.A1(_2075_),
    .A2(_2056_),
    .B1(_2023_),
    .X(_2122_));
 sky130_fd_sc_hd__or4_4 _2698_ (.A(_2119_),
    .B(_2120_),
    .C(_2121_),
    .D(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__o21a_1 _2699_ (.A1(_2002_),
    .A2(_2038_),
    .B1(_2090_),
    .X(_2124_));
 sky130_fd_sc_hd__o21a_1 _2700_ (.A1(_2088_),
    .A2(_2045_),
    .B1(_2094_),
    .X(_2125_));
 sky130_fd_sc_hd__or4_1 _2701_ (.A(_2117_),
    .B(_2123_),
    .C(_2124_),
    .D(_2125_),
    .X(_0007_));
 sky130_fd_sc_hd__buf_1 _2702_ (.A(_2008_),
    .X(_2126_));
 sky130_fd_sc_hd__or2_1 _2703_ (.A(_2101_),
    .B(_2126_),
    .X(_0008_));
 sky130_fd_sc_hd__o21a_1 _2704_ (.A1(_2106_),
    .A2(_2076_),
    .B1(_2078_),
    .X(_2127_));
 sky130_fd_sc_hd__clkbuf_2 _2705_ (.A(_2070_),
    .X(_2128_));
 sky130_fd_sc_hd__o21a_1 _2706_ (.A1(_2066_),
    .A2(_2128_),
    .B1(_2118_),
    .X(_2129_));
 sky130_fd_sc_hd__buf_1 _2707_ (.A(_2016_),
    .X(_2130_));
 sky130_fd_sc_hd__o21a_1 _2708_ (.A1(\diff3[4] ),
    .A2(_2082_),
    .B1(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__buf_1 _2709_ (.A(_2061_),
    .X(_2132_));
 sky130_fd_sc_hd__buf_1 _2710_ (.A(_2019_),
    .X(_2133_));
 sky130_fd_sc_hd__o21a_1 _2711_ (.A1(\diff3[7] ),
    .A2(_2132_),
    .B1(_2133_),
    .X(_2134_));
 sky130_fd_sc_hd__buf_1 _2712_ (.A(_2055_),
    .X(_2135_));
 sky130_fd_sc_hd__buf_1 _2713_ (.A(_2022_),
    .X(_2136_));
 sky130_fd_sc_hd__o21a_1 _2714_ (.A1(_2096_),
    .A2(_2135_),
    .B1(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__or4_4 _2715_ (.A(_2129_),
    .B(_2131_),
    .C(_2134_),
    .D(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__clkbuf_2 _2716_ (.A(_2037_),
    .X(_2139_));
 sky130_fd_sc_hd__o21a_1 _2717_ (.A1(\diff3[25] ),
    .A2(_2139_),
    .B1(_2090_),
    .X(_2140_));
 sky130_fd_sc_hd__clkbuf_2 _2718_ (.A(_2044_),
    .X(_2141_));
 sky130_fd_sc_hd__o21a_1 _2719_ (.A1(_2104_),
    .A2(_2141_),
    .B1(_2094_),
    .X(_2142_));
 sky130_fd_sc_hd__or4_4 _2720_ (.A(_2127_),
    .B(_2138_),
    .C(_2140_),
    .D(_2142_),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _2721_ (.A(_2047_),
    .B(_2126_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_1 _2722_ (.A(_2049_),
    .X(_2143_));
 sky130_fd_sc_hd__buf_1 _2723_ (.A(_2077_),
    .X(_2144_));
 sky130_fd_sc_hd__o21a_1 _2724_ (.A1(_2029_),
    .A2(_2143_),
    .B1(_2144_),
    .X(_2145_));
 sky130_fd_sc_hd__o21a_1 _2725_ (.A1(_2051_),
    .A2(_2128_),
    .B1(_2118_),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_2 _2726_ (.A(_2081_),
    .X(_2147_));
 sky130_fd_sc_hd__o21a_1 _2727_ (.A1(\diff3[5] ),
    .A2(_2147_),
    .B1(_2130_),
    .X(_2148_));
 sky130_fd_sc_hd__o21a_1 _2728_ (.A1(_2000_),
    .A2(_2132_),
    .B1(_2133_),
    .X(_2149_));
 sky130_fd_sc_hd__o21a_1 _2729_ (.A1(_2040_),
    .A2(_2135_),
    .B1(_2136_),
    .X(_2150_));
 sky130_fd_sc_hd__or4_4 _2730_ (.A(_2146_),
    .B(_2148_),
    .C(_2149_),
    .D(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__buf_1 _2731_ (.A(_2089_),
    .X(_2152_));
 sky130_fd_sc_hd__o21a_1 _2732_ (.A1(\diff3[26] ),
    .A2(_2139_),
    .B1(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__buf_1 _2733_ (.A(_2093_),
    .X(_2154_));
 sky130_fd_sc_hd__o21a_1 _2734_ (.A1(_2114_),
    .A2(_2141_),
    .B1(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__or4_4 _2735_ (.A(_2145_),
    .B(_2151_),
    .C(_2153_),
    .D(_2155_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _2736_ (.A(_2075_),
    .B(_2126_),
    .X(_0012_));
 sky130_fd_sc_hd__o21a_1 _2737_ (.A1(_2088_),
    .A2(_2143_),
    .B1(_2144_),
    .X(_2156_));
 sky130_fd_sc_hd__o21a_1 _2738_ (.A1(_2085_),
    .A2(_2128_),
    .B1(_2118_),
    .X(_2157_));
 sky130_fd_sc_hd__o21a_1 _2739_ (.A1(\diff3[6] ),
    .A2(_2147_),
    .B1(_2130_),
    .X(_2158_));
 sky130_fd_sc_hd__o21a_1 _2740_ (.A1(_2068_),
    .A2(_2132_),
    .B1(_2133_),
    .X(_2159_));
 sky130_fd_sc_hd__o21a_1 _2741_ (.A1(_2092_),
    .A2(_2135_),
    .B1(_2136_),
    .X(_2160_));
 sky130_fd_sc_hd__or4_4 _2742_ (.A(_2157_),
    .B(_2158_),
    .C(_2159_),
    .D(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__o21a_1 _2743_ (.A1(_2034_),
    .A2(_2139_),
    .B1(_2152_),
    .X(_2162_));
 sky130_fd_sc_hd__o21a_1 _2744_ (.A1(_2002_),
    .A2(_2141_),
    .B1(_2154_),
    .X(_2163_));
 sky130_fd_sc_hd__or4_4 _2745_ (.A(_2156_),
    .B(_2161_),
    .C(_2162_),
    .D(_2163_),
    .X(_0013_));
 sky130_fd_sc_hd__or2_1 _2746_ (.A(_2096_),
    .B(_2126_),
    .X(_0014_));
 sky130_fd_sc_hd__o21a_1 _2747_ (.A1(_2104_),
    .A2(_2143_),
    .B1(_2144_),
    .X(_2164_));
 sky130_fd_sc_hd__o21a_1 _2748_ (.A1(_2101_),
    .A2(_2128_),
    .B1(_2118_),
    .X(_2165_));
 sky130_fd_sc_hd__o21a_1 _2749_ (.A1(\diff3[7] ),
    .A2(_2147_),
    .B1(_2130_),
    .X(_2166_));
 sky130_fd_sc_hd__o21a_1 _2750_ (.A1(_2066_),
    .A2(_2132_),
    .B1(_2133_),
    .X(_2167_));
 sky130_fd_sc_hd__o21a_1 _2751_ (.A1(_2106_),
    .A2(_2135_),
    .B1(_2136_),
    .X(_2168_));
 sky130_fd_sc_hd__or4_4 _2752_ (.A(_2165_),
    .B(_2166_),
    .C(_2167_),
    .D(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__o21a_1 _2753_ (.A1(\diff3[28] ),
    .A2(_2139_),
    .B1(_2152_),
    .X(_2170_));
 sky130_fd_sc_hd__o21a_1 _2754_ (.A1(\diff3[25] ),
    .A2(_2141_),
    .B1(_2154_),
    .X(_2171_));
 sky130_fd_sc_hd__or4_4 _2755_ (.A(_2164_),
    .B(_2169_),
    .C(_2170_),
    .D(_2171_),
    .X(_0015_));
 sky130_fd_sc_hd__or2_1 _2756_ (.A(_2040_),
    .B(_2126_),
    .X(_0016_));
 sky130_fd_sc_hd__o21a_1 _2757_ (.A1(_2114_),
    .A2(_2143_),
    .B1(_2144_),
    .X(_2172_));
 sky130_fd_sc_hd__buf_1 _2758_ (.A(_2012_),
    .X(_2173_));
 sky130_fd_sc_hd__o21a_1 _2759_ (.A1(_2047_),
    .A2(_2128_),
    .B1(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__o21a_1 _2760_ (.A1(_2000_),
    .A2(_2147_),
    .B1(_2130_),
    .X(_2175_));
 sky130_fd_sc_hd__o21a_1 _2761_ (.A1(_2051_),
    .A2(_2132_),
    .B1(_2133_),
    .X(_2176_));
 sky130_fd_sc_hd__o21a_1 _2762_ (.A1(_2029_),
    .A2(_2135_),
    .B1(_2136_),
    .X(_2177_));
 sky130_fd_sc_hd__or4_4 _2763_ (.A(_2174_),
    .B(_2175_),
    .C(_2176_),
    .D(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__o21a_1 _2764_ (.A1(\diff3[29] ),
    .A2(_2139_),
    .B1(_2152_),
    .X(_2179_));
 sky130_fd_sc_hd__o21a_1 _2765_ (.A1(\diff3[26] ),
    .A2(_2141_),
    .B1(_2154_),
    .X(_2180_));
 sky130_fd_sc_hd__or4_4 _2766_ (.A(_2172_),
    .B(_2178_),
    .C(_2179_),
    .D(_2180_),
    .X(_0017_));
 sky130_fd_sc_hd__buf_1 _2767_ (.A(_2008_),
    .X(_2181_));
 sky130_fd_sc_hd__or2_1 _2768_ (.A(_2092_),
    .B(_2181_),
    .X(_0018_));
 sky130_fd_sc_hd__o21a_1 _2769_ (.A1(_2002_),
    .A2(_2143_),
    .B1(_2144_),
    .X(_2182_));
 sky130_fd_sc_hd__clkbuf_2 _2770_ (.A(_2070_),
    .X(_2183_));
 sky130_fd_sc_hd__o21a_1 _2771_ (.A1(_2075_),
    .A2(_2183_),
    .B1(_2173_),
    .X(_2184_));
 sky130_fd_sc_hd__buf_1 _2772_ (.A(_2016_),
    .X(_2185_));
 sky130_fd_sc_hd__o21a_1 _2773_ (.A1(_2068_),
    .A2(_2147_),
    .B1(_2185_),
    .X(_2186_));
 sky130_fd_sc_hd__clkbuf_2 _2774_ (.A(_2061_),
    .X(_2187_));
 sky130_fd_sc_hd__clkbuf_2 _2775_ (.A(_2019_),
    .X(_2188_));
 sky130_fd_sc_hd__o21a_1 _2776_ (.A1(_2085_),
    .A2(_2187_),
    .B1(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__buf_1 _2777_ (.A(_2055_),
    .X(_2190_));
 sky130_fd_sc_hd__buf_1 _2778_ (.A(_2022_),
    .X(_2191_));
 sky130_fd_sc_hd__o21a_1 _2779_ (.A1(_2088_),
    .A2(_2190_),
    .B1(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__or4_4 _2780_ (.A(_2184_),
    .B(_2186_),
    .C(_2189_),
    .D(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_2 _2781_ (.A(_2037_),
    .X(_2194_));
 sky130_fd_sc_hd__o21a_1 _2782_ (.A1(\diff3[30] ),
    .A2(_2194_),
    .B1(_2152_),
    .X(_2195_));
 sky130_fd_sc_hd__clkbuf_2 _2783_ (.A(_2044_),
    .X(_2196_));
 sky130_fd_sc_hd__o21a_1 _2784_ (.A1(_2034_),
    .A2(_2196_),
    .B1(_2154_),
    .X(_2197_));
 sky130_fd_sc_hd__or4_1 _2785_ (.A(_2182_),
    .B(_2193_),
    .C(_2195_),
    .D(_2197_),
    .X(_0019_));
 sky130_fd_sc_hd__or2_1 _2786_ (.A(_2106_),
    .B(_2181_),
    .X(_0020_));
 sky130_fd_sc_hd__buf_1 _2787_ (.A(_2049_),
    .X(_2198_));
 sky130_fd_sc_hd__buf_1 _2788_ (.A(_2077_),
    .X(_2199_));
 sky130_fd_sc_hd__o21a_1 _2789_ (.A1(\diff3[25] ),
    .A2(_2198_),
    .B1(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__o21a_1 _2790_ (.A1(_2096_),
    .A2(_2183_),
    .B1(_2173_),
    .X(_2201_));
 sky130_fd_sc_hd__clkbuf_2 _2791_ (.A(_2081_),
    .X(_2202_));
 sky130_fd_sc_hd__o21a_1 _2792_ (.A1(_2066_),
    .A2(_2202_),
    .B1(_2185_),
    .X(_2203_));
 sky130_fd_sc_hd__o21a_1 _2793_ (.A1(_2101_),
    .A2(_2187_),
    .B1(_2188_),
    .X(_2204_));
 sky130_fd_sc_hd__o21a_1 _2794_ (.A1(_2104_),
    .A2(_2190_),
    .B1(_2191_),
    .X(_2205_));
 sky130_fd_sc_hd__or4_4 _2795_ (.A(_2201_),
    .B(_2203_),
    .C(_2204_),
    .D(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__clkbuf_2 _2796_ (.A(_2089_),
    .X(_2207_));
 sky130_fd_sc_hd__o21a_1 _2797_ (.A1(\diff3[31] ),
    .A2(_2194_),
    .B1(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_2 _2798_ (.A(_2093_),
    .X(_2209_));
 sky130_fd_sc_hd__o21a_1 _2799_ (.A1(\diff3[28] ),
    .A2(_2196_),
    .B1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__or4_1 _2800_ (.A(_2200_),
    .B(_2206_),
    .C(_2208_),
    .D(_2210_),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _2801_ (.A(_2029_),
    .B(_2181_),
    .X(_0022_));
 sky130_fd_sc_hd__o21a_1 _2802_ (.A1(\diff3[26] ),
    .A2(_2198_),
    .B1(_2199_),
    .X(_2211_));
 sky130_fd_sc_hd__o21a_1 _2803_ (.A1(\diff3[17] ),
    .A2(_2183_),
    .B1(_2173_),
    .X(_2212_));
 sky130_fd_sc_hd__o21a_1 _2804_ (.A1(_2051_),
    .A2(_2202_),
    .B1(_2185_),
    .X(_2213_));
 sky130_fd_sc_hd__o21a_1 _2805_ (.A1(_2047_),
    .A2(_2187_),
    .B1(_2188_),
    .X(_2214_));
 sky130_fd_sc_hd__o21a_1 _2806_ (.A1(_2114_),
    .A2(_2190_),
    .B1(_2191_),
    .X(_2215_));
 sky130_fd_sc_hd__or4_4 _2807_ (.A(_2212_),
    .B(_2213_),
    .C(_2214_),
    .D(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__o21a_1 _2808_ (.A1(\diff3[32] ),
    .A2(_2194_),
    .B1(_2207_),
    .X(_2217_));
 sky130_fd_sc_hd__o21a_1 _2809_ (.A1(\diff3[29] ),
    .A2(_2196_),
    .B1(_2209_),
    .X(_2218_));
 sky130_fd_sc_hd__or4_4 _2810_ (.A(_2211_),
    .B(_2216_),
    .C(_2217_),
    .D(_2218_),
    .X(_0023_));
 sky130_fd_sc_hd__or2_1 _2811_ (.A(_2088_),
    .B(_2181_),
    .X(_0024_));
 sky130_fd_sc_hd__o21a_1 _2812_ (.A1(_2034_),
    .A2(_2198_),
    .B1(_2199_),
    .X(_2219_));
 sky130_fd_sc_hd__o21a_1 _2813_ (.A1(_2092_),
    .A2(_2183_),
    .B1(_2173_),
    .X(_2220_));
 sky130_fd_sc_hd__o21a_1 _2814_ (.A1(_2085_),
    .A2(_2202_),
    .B1(_2185_),
    .X(_2221_));
 sky130_fd_sc_hd__o21a_1 _2815_ (.A1(_2075_),
    .A2(_2187_),
    .B1(_2188_),
    .X(_2222_));
 sky130_fd_sc_hd__o21a_1 _2816_ (.A1(_2002_),
    .A2(_2190_),
    .B1(_2191_),
    .X(_2223_));
 sky130_fd_sc_hd__or4_4 _2817_ (.A(_2220_),
    .B(_2221_),
    .C(_2222_),
    .D(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__o21a_1 _2818_ (.A1(\diff3[33] ),
    .A2(_2194_),
    .B1(_2207_),
    .X(_2225_));
 sky130_fd_sc_hd__o21a_1 _2819_ (.A1(\diff3[30] ),
    .A2(_2196_),
    .B1(_2209_),
    .X(_2226_));
 sky130_fd_sc_hd__or4_1 _2820_ (.A(_2219_),
    .B(_2224_),
    .C(_2225_),
    .D(_2226_),
    .X(_0025_));
 sky130_fd_sc_hd__or2_1 _2821_ (.A(_2104_),
    .B(_2181_),
    .X(_0026_));
 sky130_fd_sc_hd__o21a_1 _2822_ (.A1(\diff3[28] ),
    .A2(_2198_),
    .B1(_2199_),
    .X(_2227_));
 sky130_fd_sc_hd__o21a_1 _2823_ (.A1(_2106_),
    .A2(_2183_),
    .B1(_2012_),
    .X(_2228_));
 sky130_fd_sc_hd__o21a_1 _2824_ (.A1(_2101_),
    .A2(_2202_),
    .B1(_2185_),
    .X(_2229_));
 sky130_fd_sc_hd__o21a_1 _2825_ (.A1(_2096_),
    .A2(_2187_),
    .B1(_2188_),
    .X(_2230_));
 sky130_fd_sc_hd__o21a_1 _2826_ (.A1(\diff3[25] ),
    .A2(_2190_),
    .B1(_2191_),
    .X(_2231_));
 sky130_fd_sc_hd__or4_4 _2827_ (.A(_2228_),
    .B(_2229_),
    .C(_2230_),
    .D(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__o21a_1 _2828_ (.A1(\diff3[34] ),
    .A2(_2194_),
    .B1(_2207_),
    .X(_2233_));
 sky130_fd_sc_hd__o21a_1 _2829_ (.A1(\diff3[31] ),
    .A2(_2196_),
    .B1(_2209_),
    .X(_2234_));
 sky130_fd_sc_hd__or4_1 _2830_ (.A(_2227_),
    .B(_2232_),
    .C(_2233_),
    .D(_2234_),
    .X(_0027_));
 sky130_fd_sc_hd__or2_1 _2831_ (.A(_2114_),
    .B(_2008_),
    .X(_0028_));
 sky130_fd_sc_hd__o21a_1 _2832_ (.A1(\diff3[29] ),
    .A2(_2198_),
    .B1(_2199_),
    .X(_2235_));
 sky130_fd_sc_hd__o21a_1 _2833_ (.A1(\diff3[20] ),
    .A2(_2070_),
    .B1(_2012_),
    .X(_2236_));
 sky130_fd_sc_hd__o21a_1 _2834_ (.A1(\diff3[14] ),
    .A2(_2202_),
    .B1(_2016_),
    .X(_2237_));
 sky130_fd_sc_hd__o21a_1 _2835_ (.A1(_2040_),
    .A2(_2061_),
    .B1(_2019_),
    .X(_2238_));
 sky130_fd_sc_hd__o21a_1 _2836_ (.A1(\diff3[26] ),
    .A2(_2055_),
    .B1(_2022_),
    .X(_2239_));
 sky130_fd_sc_hd__or4_4 _2837_ (.A(_2236_),
    .B(_2237_),
    .C(_2238_),
    .D(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__o21a_1 _2838_ (.A1(\diff3[35] ),
    .A2(_2037_),
    .B1(_2207_),
    .X(_2241_));
 sky130_fd_sc_hd__o21a_1 _2839_ (.A1(\diff3[32] ),
    .A2(_2044_),
    .B1(_2209_),
    .X(_2242_));
 sky130_fd_sc_hd__or4_1 _2840_ (.A(_2235_),
    .B(_2240_),
    .C(_2241_),
    .D(_2242_),
    .X(_0029_));
 sky130_fd_sc_hd__a31o_1 _2841_ (.A1(word_clk),
    .A2(_0774_),
    .A3(_0934_),
    .B1(_0031_),
    .X(_0498_));
 sky130_fd_sc_hd__inv_2 _2842_ (.A(_0000_),
    .Y(_2243_));
 sky130_fd_sc_hd__inv_2 _2843_ (.A(\word_count[14] ),
    .Y(_2244_));
 sky130_fd_sc_hd__or2_1 _2844_ (.A(net8),
    .B(net9),
    .X(_2245_));
 sky130_fd_sc_hd__or2_1 _2845_ (.A(net10),
    .B(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__or2_1 _2846_ (.A(net11),
    .B(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__or2_2 _2847_ (.A(net12),
    .B(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__or2_1 _2848_ (.A(net13),
    .B(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__or2_2 _2849_ (.A(net14),
    .B(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__or2_2 _2850_ (.A(net15),
    .B(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__or2_4 _2851_ (.A(net16),
    .B(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__or3_1 _2852_ (.A(net2),
    .B(net3),
    .C(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__or2_2 _2853_ (.A(net4),
    .B(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__or2_1 _2854_ (.A(net5),
    .B(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__or2_2 _2855_ (.A(net6),
    .B(_2255_),
    .X(_2256_));
 sky130_fd_sc_hd__or4_4 _2856_ (.A(net6),
    .B(net7),
    .C(net4),
    .D(net5),
    .X(_2257_));
 sky130_fd_sc_hd__buf_1 _2857_ (.A(_2253_),
    .X(_2258_));
 sky130_fd_sc_hd__or2_2 _2858_ (.A(_2257_),
    .B(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__inv_2 _2859_ (.A(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__a21oi_2 _2860_ (.A1(net7),
    .A2(_2256_),
    .B1(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__inv_2 _2861_ (.A(_2261_),
    .Y(_2262_));
 sky130_fd_sc_hd__o22a_1 _2862_ (.A1(_2244_),
    .A2(_2261_),
    .B1(\word_count[14] ),
    .B2(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__a21boi_2 _2863_ (.A1(net5),
    .A2(_2254_),
    .B1_N(_2255_),
    .Y(_2264_));
 sky130_fd_sc_hd__inv_2 _2864_ (.A(net3),
    .Y(_2265_));
 sky130_fd_sc_hd__buf_2 _2865_ (.A(net2),
    .X(_2266_));
 sky130_fd_sc_hd__nor2_4 _2866_ (.A(_2266_),
    .B(_2252_),
    .Y(_2267_));
 sky130_fd_sc_hd__o21ai_1 _2867_ (.A1(_2265_),
    .A2(_2267_),
    .B1(_2258_),
    .Y(_2268_));
 sky130_fd_sc_hd__o2bb2a_1 _2868_ (.A1_N(\word_count[10] ),
    .A2_N(_2268_),
    .B1(\word_count[10] ),
    .B2(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__clkbuf_2 _2869_ (.A(\word_count[9] ),
    .X(_2270_));
 sky130_fd_sc_hd__a21oi_4 _2870_ (.A1(_2266_),
    .A2(_2252_),
    .B1(_2267_),
    .Y(_2271_));
 sky130_fd_sc_hd__clkbuf_2 _2871_ (.A(\word_count[8] ),
    .X(_2272_));
 sky130_fd_sc_hd__a21boi_2 _2872_ (.A1(net16),
    .A2(_2251_),
    .B1_N(_2252_),
    .Y(_2273_));
 sky130_fd_sc_hd__a22oi_2 _2873_ (.A1(_2272_),
    .A2(_2273_),
    .B1(_2270_),
    .B2(_2271_),
    .Y(_2274_));
 sky130_fd_sc_hd__o221ai_2 _2874_ (.A1(_2270_),
    .A2(_2271_),
    .B1(\word_count[12] ),
    .B2(_2264_),
    .C1(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__inv_2 _2875_ (.A(\word_count[13] ),
    .Y(_2276_));
 sky130_fd_sc_hd__a21bo_1 _2876_ (.A1(net6),
    .A2(_2255_),
    .B1_N(_2256_),
    .X(_2277_));
 sky130_fd_sc_hd__inv_2 _2877_ (.A(\word_count[11] ),
    .Y(_2278_));
 sky130_fd_sc_hd__a21bo_1 _2878_ (.A1(net4),
    .A2(_2258_),
    .B1_N(_2254_),
    .X(_2279_));
 sky130_fd_sc_hd__inv_2 _2879_ (.A(_2279_),
    .Y(_2280_));
 sky130_fd_sc_hd__inv_2 _2880_ (.A(\word_count[15] ),
    .Y(_2281_));
 sky130_fd_sc_hd__inv_2 _2881_ (.A(net14),
    .Y(_2282_));
 sky130_fd_sc_hd__inv_2 _2882_ (.A(_2249_),
    .Y(_2283_));
 sky130_fd_sc_hd__o21ai_2 _2883_ (.A1(_2282_),
    .A2(_2283_),
    .B1(_2250_),
    .Y(_2284_));
 sky130_fd_sc_hd__inv_2 _2884_ (.A(\word_count[6] ),
    .Y(_2285_));
 sky130_fd_sc_hd__inv_2 _2885_ (.A(_2284_),
    .Y(_2286_));
 sky130_fd_sc_hd__a22o_1 _2886_ (.A1(\word_count[6] ),
    .A2(_2284_),
    .B1(_2285_),
    .B2(_2286_),
    .X(_2287_));
 sky130_fd_sc_hd__o221a_1 _2887_ (.A1(\word_count[15] ),
    .A2(_2259_),
    .B1(_2281_),
    .B2(_2260_),
    .C1(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__a21bo_1 _2888_ (.A1(net15),
    .A2(_2250_),
    .B1_N(_2251_),
    .X(_2289_));
 sky130_fd_sc_hd__inv_2 _2889_ (.A(_2289_),
    .Y(_2290_));
 sky130_fd_sc_hd__inv_2 _2890_ (.A(\word_count[7] ),
    .Y(_2291_));
 sky130_fd_sc_hd__clkbuf_2 _2891_ (.A(net13),
    .X(_2292_));
 sky130_fd_sc_hd__a21oi_4 _2892_ (.A1(_2292_),
    .A2(_2248_),
    .B1(_2283_),
    .Y(_2293_));
 sky130_fd_sc_hd__inv_2 _2893_ (.A(\word_count[5] ),
    .Y(_2294_));
 sky130_fd_sc_hd__inv_2 _2894_ (.A(_2293_),
    .Y(_2295_));
 sky130_fd_sc_hd__inv_2 _2895_ (.A(\word_count[2] ),
    .Y(_2296_));
 sky130_fd_sc_hd__a21bo_1 _2896_ (.A1(net10),
    .A2(_2245_),
    .B1_N(_2246_),
    .X(_2297_));
 sky130_fd_sc_hd__inv_2 _2897_ (.A(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__inv_2 _2898_ (.A(\word_count[0] ),
    .Y(_2299_));
 sky130_fd_sc_hd__buf_1 _2899_ (.A(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__inv_2 _2900_ (.A(\word_count[1] ),
    .Y(_2301_));
 sky130_fd_sc_hd__a2bb2o_1 _2901_ (.A1_N(_2301_),
    .A2_N(net9),
    .B1(_2301_),
    .B2(net9),
    .X(_2302_));
 sky130_fd_sc_hd__inv_2 _2902_ (.A(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__nand2_1 _2903_ (.A(_2299_),
    .B(net8),
    .Y(_2304_));
 sky130_fd_sc_hd__o32a_1 _2904_ (.A1(_2300_),
    .A2(net8),
    .A3(_2303_),
    .B1(_2302_),
    .B2(_2304_),
    .X(_2305_));
 sky130_fd_sc_hd__a221o_1 _2905_ (.A1(_2296_),
    .A2(_2297_),
    .B1(\word_count[2] ),
    .B2(_2298_),
    .C1(_2305_),
    .X(_2306_));
 sky130_fd_sc_hd__buf_1 _2906_ (.A(\word_count[3] ),
    .X(_2307_));
 sky130_fd_sc_hd__inv_2 _2907_ (.A(_2247_),
    .Y(_2308_));
 sky130_fd_sc_hd__a21o_1 _2908_ (.A1(net11),
    .A2(_2246_),
    .B1(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__o2bb2a_1 _2909_ (.A1_N(_2307_),
    .A2_N(_2309_),
    .B1(_2307_),
    .B2(_2309_),
    .X(_2310_));
 sky130_fd_sc_hd__buf_1 _2910_ (.A(\word_count[4] ),
    .X(_2311_));
 sky130_fd_sc_hd__inv_2 _2911_ (.A(net12),
    .Y(_2312_));
 sky130_fd_sc_hd__o21ai_1 _2912_ (.A1(_2312_),
    .A2(_2308_),
    .B1(_2248_),
    .Y(_2313_));
 sky130_fd_sc_hd__o2bb2a_1 _2913_ (.A1_N(_2311_),
    .A2_N(_2313_),
    .B1(_2311_),
    .B2(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__or3_1 _2914_ (.A(_2306_),
    .B(_2310_),
    .C(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__a221oi_2 _2915_ (.A1(\word_count[5] ),
    .A2(_2293_),
    .B1(_2294_),
    .B2(_2295_),
    .C1(_2315_),
    .Y(_2316_));
 sky130_fd_sc_hd__o221a_1 _2916_ (.A1(\word_count[7] ),
    .A2(_2290_),
    .B1(_2291_),
    .B2(_2289_),
    .C1(_2316_),
    .X(_2317_));
 sky130_fd_sc_hd__o211a_1 _2917_ (.A1(_2272_),
    .A2(_2273_),
    .B1(_2288_),
    .C1(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__o221a_1 _2918_ (.A1(_2278_),
    .A2(_2279_),
    .B1(\word_count[11] ),
    .B2(_2280_),
    .C1(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__o21ai_1 _2919_ (.A1(_2276_),
    .A2(_2277_),
    .B1(_2319_),
    .Y(_2320_));
 sky130_fd_sc_hd__a21o_1 _2920_ (.A1(_2276_),
    .A2(_2277_),
    .B1(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__a2111o_4 _2921_ (.A1(\word_count[12] ),
    .A2(_2264_),
    .B1(_2269_),
    .C1(_2275_),
    .D1(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__nor3_4 _2922_ (.A(_2263_),
    .B(_2322_),
    .C(_2260_),
    .Y(_0031_));
 sky130_fd_sc_hd__nand2_1 _2923_ (.A(enable),
    .B(_0031_),
    .Y(_2323_));
 sky130_fd_sc_hd__clkbuf_4 _2924_ (.A(net18),
    .X(_2324_));
 sky130_fd_sc_hd__a221o_1 _2925_ (.A1(enable),
    .A2(_2243_),
    .B1(_0000_),
    .B2(_2323_),
    .C1(_2324_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_mclk1 (.A(mclk1),
    .X(clknet_0_mclk1));
 sky130_fd_sc_hd__buf_1 _2927_ (.A(net41),
    .X(_2326_));
 sky130_fd_sc_hd__buf_1 _2928_ (.A(_2326_),
    .X(_0146_));
 sky130_fd_sc_hd__clkinvlp_2 _2929_ (.A(\acc1[36] ),
    .Y(_2327_));
 sky130_fd_sc_hd__inv_2 _2930_ (.A(\acc2[36] ),
    .Y(_2328_));
 sky130_fd_sc_hd__o22a_1 _2931_ (.A1(\acc1[36] ),
    .A2(\acc2[36] ),
    .B1(_2327_),
    .B2(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__nor2_1 _2932_ (.A(\acc1[35] ),
    .B(\acc2[35] ),
    .Y(_2330_));
 sky130_fd_sc_hd__a21oi_2 _2933_ (.A1(\acc1[35] ),
    .A2(\acc2[35] ),
    .B1(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__inv_2 _2934_ (.A(_2331_),
    .Y(_2332_));
 sky130_fd_sc_hd__clkinvlp_4 _2935_ (.A(\acc1[34] ),
    .Y(_2333_));
 sky130_fd_sc_hd__inv_2 _2936_ (.A(\acc2[34] ),
    .Y(_2334_));
 sky130_fd_sc_hd__clkbuf_2 _2937_ (.A(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__o22a_1 _2938_ (.A1(_2333_),
    .A2(_2335_),
    .B1(\acc1[34] ),
    .B2(\acc2[34] ),
    .X(_2336_));
 sky130_fd_sc_hd__inv_2 _2939_ (.A(_2336_),
    .Y(_2337_));
 sky130_fd_sc_hd__nor2_1 _2940_ (.A(\acc1[33] ),
    .B(\acc2[33] ),
    .Y(_2338_));
 sky130_fd_sc_hd__a21oi_2 _2941_ (.A1(\acc1[33] ),
    .A2(\acc2[33] ),
    .B1(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__inv_2 _2942_ (.A(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__clkinvlp_4 _2943_ (.A(\acc1[32] ),
    .Y(_2341_));
 sky130_fd_sc_hd__inv_2 _2944_ (.A(\acc2[32] ),
    .Y(_2342_));
 sky130_fd_sc_hd__clkbuf_2 _2945_ (.A(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__o22a_1 _2946_ (.A1(_2341_),
    .A2(_2343_),
    .B1(\acc1[32] ),
    .B2(\acc2[32] ),
    .X(_2344_));
 sky130_fd_sc_hd__inv_2 _2947_ (.A(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__clkinv_1 _2948_ (.A(\acc1[28] ),
    .Y(_2346_));
 sky130_fd_sc_hd__inv_2 _2949_ (.A(\acc2[28] ),
    .Y(_2347_));
 sky130_fd_sc_hd__o22a_1 _2950_ (.A1(\acc1[28] ),
    .A2(\acc2[28] ),
    .B1(_2346_),
    .B2(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__inv_2 _2951_ (.A(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__clkbuf_2 _2952_ (.A(\acc2[29] ),
    .X(_2350_));
 sky130_fd_sc_hd__clkinv_1 _2953_ (.A(\acc1[29] ),
    .Y(_2351_));
 sky130_fd_sc_hd__inv_2 _2954_ (.A(\acc2[29] ),
    .Y(_2352_));
 sky130_fd_sc_hd__o22a_1 _2955_ (.A1(\acc1[29] ),
    .A2(_2350_),
    .B1(_2351_),
    .B2(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__inv_2 _2956_ (.A(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__or2_1 _2957_ (.A(_2349_),
    .B(_2354_),
    .X(_2355_));
 sky130_fd_sc_hd__clkinvlp_4 _2958_ (.A(\acc1[30] ),
    .Y(_2356_));
 sky130_fd_sc_hd__inv_2 _2959_ (.A(\acc2[30] ),
    .Y(_2357_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2960_ (.A(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__o22a_1 _2961_ (.A1(\acc1[30] ),
    .A2(\acc2[30] ),
    .B1(_2356_),
    .B2(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__nor2_1 _2962_ (.A(\acc1[31] ),
    .B(\acc2[31] ),
    .Y(_2360_));
 sky130_fd_sc_hd__a21oi_2 _2963_ (.A1(\acc1[31] ),
    .A2(\acc2[31] ),
    .B1(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__nand2_1 _2964_ (.A(_2359_),
    .B(_2361_),
    .Y(_2362_));
 sky130_fd_sc_hd__or2_1 _2965_ (.A(_2355_),
    .B(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__inv_1 _2966_ (.A(\acc1[27] ),
    .Y(_2364_));
 sky130_fd_sc_hd__inv_2 _2967_ (.A(\acc2[27] ),
    .Y(_2365_));
 sky130_fd_sc_hd__clkbuf_2 _2968_ (.A(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__o22a_1 _2969_ (.A1(_2364_),
    .A2(_2366_),
    .B1(\acc1[27] ),
    .B2(\acc2[27] ),
    .X(_2367_));
 sky130_fd_sc_hd__inv_6 _2970_ (.A(\acc1[26] ),
    .Y(_2368_));
 sky130_fd_sc_hd__inv_2 _2971_ (.A(\acc2[26] ),
    .Y(_2369_));
 sky130_fd_sc_hd__clkbuf_2 _2972_ (.A(_2369_),
    .X(_0499_));
 sky130_fd_sc_hd__o22a_1 _2973_ (.A1(_2368_),
    .A2(_0499_),
    .B1(\acc1[26] ),
    .B2(\acc2[26] ),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _2974_ (.A(_2367_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__clkinv_1 _2975_ (.A(\acc1[25] ),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _2976_ (.A(\acc2[25] ),
    .Y(_0503_));
 sky130_fd_sc_hd__clkbuf_2 _2977_ (.A(\acc2[25] ),
    .X(_0504_));
 sky130_fd_sc_hd__o22a_1 _2978_ (.A1(_0502_),
    .A2(_0503_),
    .B1(\acc1[25] ),
    .B2(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__inv_2 _2979_ (.A(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__clkinv_1 _2980_ (.A(\acc1[24] ),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_2 _2981_ (.A(\acc2[24] ),
    .Y(_0508_));
 sky130_fd_sc_hd__o22a_1 _2982_ (.A1(_0507_),
    .A2(_0508_),
    .B1(\acc1[24] ),
    .B2(\acc2[24] ),
    .X(_0509_));
 sky130_fd_sc_hd__inv_2 _2983_ (.A(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__or2_1 _2984_ (.A(_0506_),
    .B(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__or2_1 _2985_ (.A(_0501_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_2 _2986_ (.A(\acc1[23] ),
    .B(\acc2[23] ),
    .Y(_0513_));
 sky130_fd_sc_hd__clkinv_1 _2987_ (.A(\acc1[23] ),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_2 _2988_ (.A(\acc2[23] ),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_1 _2989_ (.A(\acc1[22] ),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _2990_ (.A(\acc2[22] ),
    .Y(_0517_));
 sky130_fd_sc_hd__clkbuf_2 _2991_ (.A(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_2 _2992_ (.A(\acc2[21] ),
    .X(_0519_));
 sky130_fd_sc_hd__clkinv_1 _2993_ (.A(\acc1[21] ),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _2994_ (.A(\acc2[21] ),
    .Y(_0521_));
 sky130_fd_sc_hd__o22a_1 _2995_ (.A1(\acc1[21] ),
    .A2(_0519_),
    .B1(_0520_),
    .B2(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__inv_2 _2996_ (.A(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__clkinv_1 _2997_ (.A(\acc1[20] ),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _2998_ (.A(\acc2[20] ),
    .Y(_0525_));
 sky130_fd_sc_hd__o22a_1 _2999_ (.A1(_0524_),
    .A2(_0525_),
    .B1(\acc1[20] ),
    .B2(\acc2[20] ),
    .X(_0526_));
 sky130_fd_sc_hd__inv_2 _3000_ (.A(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__or2_1 _3001_ (.A(_0523_),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__inv_1 _3002_ (.A(\acc1[19] ),
    .Y(_0529_));
 sky130_fd_sc_hd__inv_2 _3003_ (.A(\acc2[19] ),
    .Y(_0530_));
 sky130_fd_sc_hd__clkbuf_2 _3004_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__o22a_1 _3005_ (.A1(\acc1[19] ),
    .A2(\acc2[19] ),
    .B1(_0529_),
    .B2(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__clkinvlp_4 _3006_ (.A(\acc1[18] ),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _3007_ (.A(\acc2[18] ),
    .Y(_0534_));
 sky130_fd_sc_hd__clkbuf_2 _3008_ (.A(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__o22a_1 _3009_ (.A1(_0533_),
    .A2(_0535_),
    .B1(\acc1[18] ),
    .B2(\acc2[18] ),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _3010_ (.A(_0532_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__clkbuf_2 _3011_ (.A(\acc2[17] ),
    .X(_0538_));
 sky130_fd_sc_hd__a22o_1 _3012_ (.A1(\acc1[17] ),
    .A2(_0538_),
    .B1(\acc1[16] ),
    .B2(\acc2[16] ),
    .X(_0539_));
 sky130_fd_sc_hd__o21ai_1 _3013_ (.A1(\acc1[17] ),
    .A2(_0538_),
    .B1(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__a211o_1 _3014_ (.A1(_0529_),
    .A2(_0531_),
    .B1(_0533_),
    .C1(_0535_),
    .X(_0541_));
 sky130_fd_sc_hd__o221a_1 _3015_ (.A1(_0529_),
    .A2(_0531_),
    .B1(_0537_),
    .B2(_0540_),
    .C1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__or2_1 _3016_ (.A(_0528_),
    .B(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _3017_ (.A1(\acc1[21] ),
    .A2(_0519_),
    .B1(\acc1[20] ),
    .B2(\acc2[20] ),
    .X(_0544_));
 sky130_fd_sc_hd__o21ai_1 _3018_ (.A1(\acc1[21] ),
    .A2(_0519_),
    .B1(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a22o_1 _3019_ (.A1(_0516_),
    .A2(_0518_),
    .B1(_0543_),
    .B2(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__o221a_1 _3020_ (.A1(_0514_),
    .A2(_0515_),
    .B1(_0516_),
    .B2(_0518_),
    .C1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_1 _3021_ (.A(\acc1[15] ),
    .B(\acc2[15] ),
    .Y(_0548_));
 sky130_fd_sc_hd__a21oi_2 _3022_ (.A1(\acc1[15] ),
    .A2(\acc2[15] ),
    .B1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__clkinvlp_4 _3023_ (.A(\acc1[14] ),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_2 _3024_ (.A(\acc2[14] ),
    .Y(_0551_));
 sky130_fd_sc_hd__clkbuf_2 _3025_ (.A(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__o22a_1 _3026_ (.A1(_0550_),
    .A2(_0552_),
    .B1(\acc1[14] ),
    .B2(\acc2[14] ),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_1 _3027_ (.A(_0549_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__clkinv_1 _3028_ (.A(\acc1[13] ),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_2 _3029_ (.A(\acc2[13] ),
    .Y(_0556_));
 sky130_fd_sc_hd__clkbuf_2 _3030_ (.A(\acc2[13] ),
    .X(_0557_));
 sky130_fd_sc_hd__o22a_1 _3031_ (.A1(_0555_),
    .A2(_0556_),
    .B1(\acc1[13] ),
    .B2(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__inv_2 _3032_ (.A(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__clkinv_1 _3033_ (.A(\acc1[12] ),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_2 _3034_ (.A(\acc2[12] ),
    .Y(_0561_));
 sky130_fd_sc_hd__o22a_1 _3035_ (.A1(_0560_),
    .A2(_0561_),
    .B1(\acc1[12] ),
    .B2(\acc2[12] ),
    .X(_0562_));
 sky130_fd_sc_hd__inv_2 _3036_ (.A(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__or2_1 _3037_ (.A(_0559_),
    .B(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__or2_1 _3038_ (.A(_0554_),
    .B(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__inv_1 _3039_ (.A(\acc1[11] ),
    .Y(_0566_));
 sky130_fd_sc_hd__inv_2 _3040_ (.A(\acc2[11] ),
    .Y(_0567_));
 sky130_fd_sc_hd__clkbuf_2 _3041_ (.A(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__o22a_1 _3042_ (.A1(_0566_),
    .A2(_0568_),
    .B1(\acc1[11] ),
    .B2(\acc2[11] ),
    .X(_0569_));
 sky130_fd_sc_hd__clkinvlp_4 _3043_ (.A(\acc1[10] ),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_2 _3044_ (.A(\acc2[10] ),
    .Y(_0571_));
 sky130_fd_sc_hd__clkbuf_2 _3045_ (.A(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__o22a_1 _3046_ (.A1(_0570_),
    .A2(_0572_),
    .B1(\acc1[10] ),
    .B2(\acc2[10] ),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_1 _3047_ (.A(_0569_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__clkinv_1 _3048_ (.A(\acc1[9] ),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_2 _3049_ (.A(\acc2[9] ),
    .Y(_0576_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3050_ (.A(\acc2[9] ),
    .X(_0577_));
 sky130_fd_sc_hd__o22a_1 _3051_ (.A1(_0575_),
    .A2(_0576_),
    .B1(\acc1[9] ),
    .B2(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__inv_2 _3052_ (.A(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__clkinv_1 _3053_ (.A(\acc1[8] ),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_2 _3054_ (.A(\acc2[8] ),
    .Y(_0581_));
 sky130_fd_sc_hd__o22a_1 _3055_ (.A1(_0580_),
    .A2(_0581_),
    .B1(\acc1[8] ),
    .B2(\acc2[8] ),
    .X(_0582_));
 sky130_fd_sc_hd__inv_2 _3056_ (.A(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__or2_1 _3057_ (.A(_0579_),
    .B(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__or2_1 _3058_ (.A(_0574_),
    .B(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__nor2_1 _3059_ (.A(\acc1[7] ),
    .B(\acc2[7] ),
    .Y(_0586_));
 sky130_fd_sc_hd__a21oi_2 _3060_ (.A1(\acc1[7] ),
    .A2(\acc2[7] ),
    .B1(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__inv_2 _3061_ (.A(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__clkinvlp_4 _3062_ (.A(\acc1[6] ),
    .Y(_0589_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(\acc2[6] ),
    .Y(_0590_));
 sky130_fd_sc_hd__clkbuf_2 _3064_ (.A(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__o22a_1 _3065_ (.A1(_0589_),
    .A2(_0591_),
    .B1(\acc1[6] ),
    .B2(\acc2[6] ),
    .X(_0592_));
 sky130_fd_sc_hd__inv_2 _3066_ (.A(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(\acc1[5] ),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_2 _3068_ (.A(\acc2[5] ),
    .Y(_0595_));
 sky130_fd_sc_hd__nor2_2 _3069_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _3070_ (.A(\acc1[4] ),
    .Y(_0597_));
 sky130_fd_sc_hd__clkinv_4 _3071_ (.A(\acc2[4] ),
    .Y(_0598_));
 sky130_fd_sc_hd__nor2_4 _3072_ (.A(_0597_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__o22a_1 _3073_ (.A1(\acc1[5] ),
    .A2(\acc2[5] ),
    .B1(_0596_),
    .B2(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__clkinv_1 _3075_ (.A(\acc1[7] ),
    .Y(_0602_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(\acc2[7] ),
    .Y(_0603_));
 sky130_fd_sc_hd__o32a_1 _3077_ (.A1(_0589_),
    .A2(_0591_),
    .A3(_0586_),
    .B1(_0602_),
    .B2(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__a21oi_4 _3078_ (.A1(_0594_),
    .A2(_0595_),
    .B1(_0596_),
    .Y(_0605_));
 sky130_fd_sc_hd__a21oi_4 _3079_ (.A1(_0597_),
    .A2(_0598_),
    .B1(_0599_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _3080_ (.A(_0605_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor2_1 _3081_ (.A(\acc1[3] ),
    .B(\acc2[3] ),
    .Y(_0608_));
 sky130_fd_sc_hd__a21oi_2 _3082_ (.A1(\acc1[3] ),
    .A2(\acc2[3] ),
    .B1(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__inv_2 _3083_ (.A(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__inv_1 _3084_ (.A(\acc1[2] ),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _3085_ (.A(\acc2[2] ),
    .Y(_0612_));
 sky130_fd_sc_hd__clkbuf_2 _3086_ (.A(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__o22a_1 _3087_ (.A1(_0611_),
    .A2(_0613_),
    .B1(\acc1[2] ),
    .B2(\acc2[2] ),
    .X(_0614_));
 sky130_fd_sc_hd__inv_2 _3088_ (.A(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__clkinvlp_2 _3089_ (.A(\acc1[1] ),
    .Y(_0616_));
 sky130_fd_sc_hd__clkbuf_2 _3090_ (.A(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _3091_ (.A(\acc2[1] ),
    .Y(_0618_));
 sky130_fd_sc_hd__clkinv_1 _3092_ (.A(\acc1[0] ),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_2 _3093_ (.A(\acc2[0] ),
    .Y(_0620_));
 sky130_fd_sc_hd__clkbuf_2 _3094_ (.A(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__a22o_1 _3095_ (.A1(\acc1[1] ),
    .A2(\acc2[1] ),
    .B1(_0617_),
    .B2(_0618_),
    .X(_0622_));
 sky130_fd_sc_hd__or3_1 _3096_ (.A(_0619_),
    .B(_0621_),
    .C(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__o21ai_2 _3097_ (.A1(_0617_),
    .A2(_0618_),
    .B1(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__inv_2 _3098_ (.A(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__clkinvlp_2 _3099_ (.A(\acc1[3] ),
    .Y(_0626_));
 sky130_fd_sc_hd__inv_2 _3100_ (.A(\acc2[3] ),
    .Y(_0627_));
 sky130_fd_sc_hd__o32a_1 _3101_ (.A1(_0611_),
    .A2(_0613_),
    .A3(_0608_),
    .B1(_0626_),
    .B2(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__o31a_1 _3102_ (.A1(_0610_),
    .A2(_0615_),
    .A3(_0625_),
    .B1(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__or4_4 _3103_ (.A(_0588_),
    .B(_0593_),
    .C(_0607_),
    .D(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__o311a_2 _3104_ (.A1(_0588_),
    .A2(_0593_),
    .A3(_0601_),
    .B1(_0604_),
    .C1(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__a22o_1 _3105_ (.A1(\acc1[13] ),
    .A2(_0557_),
    .B1(\acc1[12] ),
    .B2(\acc2[12] ),
    .X(_0632_));
 sky130_fd_sc_hd__o21ai_1 _3106_ (.A1(\acc1[13] ),
    .A2(_0557_),
    .B1(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__a22o_1 _3107_ (.A1(\acc1[9] ),
    .A2(_0577_),
    .B1(\acc1[8] ),
    .B2(\acc2[8] ),
    .X(_0634_));
 sky130_fd_sc_hd__o21ai_1 _3108_ (.A1(\acc1[9] ),
    .A2(_0577_),
    .B1(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__a211o_1 _3109_ (.A1(_0566_),
    .A2(_0568_),
    .B1(_0570_),
    .C1(_0572_),
    .X(_0636_));
 sky130_fd_sc_hd__o221a_1 _3110_ (.A1(_0566_),
    .A2(_0568_),
    .B1(_0574_),
    .B2(_0635_),
    .C1(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__inv_2 _3111_ (.A(\acc1[15] ),
    .Y(_0638_));
 sky130_fd_sc_hd__inv_2 _3112_ (.A(\acc2[15] ),
    .Y(_0639_));
 sky130_fd_sc_hd__o32a_1 _3113_ (.A1(_0550_),
    .A2(_0552_),
    .A3(_0548_),
    .B1(_0638_),
    .B2(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__o221a_1 _3114_ (.A1(_0554_),
    .A2(_0633_),
    .B1(_0565_),
    .B2(_0637_),
    .C1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__o31a_2 _3115_ (.A1(_0565_),
    .A2(_0585_),
    .A3(_0631_),
    .B1(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__inv_2 _3116_ (.A(\acc1[17] ),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_2 _3117_ (.A(\acc2[17] ),
    .Y(_0644_));
 sky130_fd_sc_hd__o22a_1 _3118_ (.A1(\acc1[17] ),
    .A2(_0538_),
    .B1(_0643_),
    .B2(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__inv_2 _3119_ (.A(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__clkinv_1 _3120_ (.A(\acc1[16] ),
    .Y(_0647_));
 sky130_fd_sc_hd__inv_2 _3121_ (.A(\acc2[16] ),
    .Y(_0648_));
 sky130_fd_sc_hd__o22a_1 _3122_ (.A1(_0647_),
    .A2(_0648_),
    .B1(\acc1[16] ),
    .B2(\acc2[16] ),
    .X(_0649_));
 sky130_fd_sc_hd__inv_2 _3123_ (.A(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__or2_1 _3124_ (.A(_0646_),
    .B(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__or2_1 _3125_ (.A(_0537_),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__a21oi_2 _3126_ (.A1(\acc1[23] ),
    .A2(\acc2[23] ),
    .B1(_0513_),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_2 _3127_ (.A(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__o22a_1 _3128_ (.A1(\acc1[22] ),
    .A2(\acc2[22] ),
    .B1(_0516_),
    .B2(_0517_),
    .X(_0655_));
 sky130_fd_sc_hd__or4b_4 _3129_ (.A(_0652_),
    .B(_0654_),
    .C(_0528_),
    .D_N(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__o22a_2 _3130_ (.A1(_0513_),
    .A2(_0547_),
    .B1(_0642_),
    .B2(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__a22o_1 _3131_ (.A1(\acc1[28] ),
    .A2(\acc2[28] ),
    .B1(\acc1[29] ),
    .B2(_2350_),
    .X(_0658_));
 sky130_fd_sc_hd__o21ai_1 _3132_ (.A1(\acc1[29] ),
    .A2(_2350_),
    .B1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__a22o_1 _3133_ (.A1(\acc1[25] ),
    .A2(_0504_),
    .B1(\acc1[24] ),
    .B2(\acc2[24] ),
    .X(_0660_));
 sky130_fd_sc_hd__o21ai_1 _3134_ (.A1(\acc1[25] ),
    .A2(_0504_),
    .B1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__a211o_1 _3135_ (.A1(_2364_),
    .A2(_2366_),
    .B1(_2368_),
    .C1(_0499_),
    .X(_0662_));
 sky130_fd_sc_hd__o221a_1 _3136_ (.A1(_2364_),
    .A2(_2366_),
    .B1(_0501_),
    .B2(_0661_),
    .C1(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__clkinv_1 _3137_ (.A(\acc1[31] ),
    .Y(_0664_));
 sky130_fd_sc_hd__inv_2 _3138_ (.A(\acc2[31] ),
    .Y(_0665_));
 sky130_fd_sc_hd__o32a_1 _3139_ (.A1(_2356_),
    .A2(_2358_),
    .A3(_2360_),
    .B1(_0664_),
    .B2(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__o221a_1 _3140_ (.A1(_2362_),
    .A2(_0659_),
    .B1(_2363_),
    .B2(_0663_),
    .C1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__o31a_1 _3141_ (.A1(_2363_),
    .A2(_0512_),
    .A3(_0657_),
    .B1(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__clkinv_1 _3142_ (.A(\acc1[33] ),
    .Y(_0669_));
 sky130_fd_sc_hd__inv_2 _3143_ (.A(\acc2[33] ),
    .Y(_0670_));
 sky130_fd_sc_hd__o32a_1 _3144_ (.A1(_2341_),
    .A2(_2343_),
    .A3(_2338_),
    .B1(_0669_),
    .B2(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__o31a_1 _3145_ (.A1(_2340_),
    .A2(_2345_),
    .A3(_0668_),
    .B1(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__inv_2 _3146_ (.A(\acc1[35] ),
    .Y(_0673_));
 sky130_fd_sc_hd__inv_2 _3147_ (.A(\acc2[35] ),
    .Y(_0674_));
 sky130_fd_sc_hd__o32a_1 _3148_ (.A1(_2333_),
    .A2(_2335_),
    .A3(_2330_),
    .B1(_0673_),
    .B2(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__o31a_1 _3149_ (.A1(_2332_),
    .A2(_2337_),
    .A3(_0672_),
    .B1(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__inv_2 _3150_ (.A(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_2 _3151_ (.A(_2329_),
    .Y(_0678_));
 sky130_fd_sc_hd__inv_2 _3152_ (.A(net18),
    .Y(_0679_));
 sky130_fd_sc_hd__clkbuf_2 _3153_ (.A(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_2 _3154_ (.A(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_2 _3155_ (.A(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__o221a_1 _3156_ (.A1(_2329_),
    .A2(_0677_),
    .B1(_0678_),
    .B2(_0676_),
    .C1(_0682_),
    .X(_0496_));
 sky130_fd_sc_hd__buf_1 _3157_ (.A(_0146_),
    .X(_0145_));
 sky130_fd_sc_hd__or2_1 _3158_ (.A(_0672_),
    .B(_2337_),
    .X(_0683_));
 sky130_fd_sc_hd__o21ai_1 _3159_ (.A1(_2333_),
    .A2(_2335_),
    .B1(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _3160_ (.A(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__o221a_1 _3161_ (.A1(_2332_),
    .A2(_0685_),
    .B1(_2331_),
    .B2(_0684_),
    .C1(_0682_),
    .X(_0495_));
 sky130_fd_sc_hd__buf_1 _3162_ (.A(_0146_),
    .X(_0144_));
 sky130_fd_sc_hd__inv_2 _3163_ (.A(_0672_),
    .Y(_0686_));
 sky130_fd_sc_hd__clkbuf_2 _3164_ (.A(_0679_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_4 _3165_ (.A(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__o211a_1 _3166_ (.A1(_0686_),
    .A2(_2336_),
    .B1(_0688_),
    .C1(_0683_),
    .X(_0494_));
 sky130_fd_sc_hd__buf_1 _3167_ (.A(_0146_),
    .X(_0143_));
 sky130_fd_sc_hd__or2_1 _3168_ (.A(_0668_),
    .B(_2345_),
    .X(_0689_));
 sky130_fd_sc_hd__o21ai_1 _3169_ (.A1(_2341_),
    .A2(_2343_),
    .B1(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__inv_2 _3170_ (.A(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__o221a_1 _3171_ (.A1(_2340_),
    .A2(_0691_),
    .B1(_2339_),
    .B2(_0690_),
    .C1(_0682_),
    .X(_0493_));
 sky130_fd_sc_hd__buf_1 _3172_ (.A(_0146_),
    .X(_0142_));
 sky130_fd_sc_hd__inv_2 _3173_ (.A(_0668_),
    .Y(_0692_));
 sky130_fd_sc_hd__o211a_1 _3174_ (.A1(_0692_),
    .A2(_2344_),
    .B1(_0688_),
    .C1(_0689_),
    .X(_0492_));
 sky130_fd_sc_hd__buf_1 _3175_ (.A(_2326_),
    .X(_0693_));
 sky130_fd_sc_hd__buf_1 _3176_ (.A(_0693_),
    .X(_0141_));
 sky130_fd_sc_hd__o21ai_1 _3177_ (.A1(_0657_),
    .A2(_0512_),
    .B1(_0663_),
    .Y(_0694_));
 sky130_fd_sc_hd__inv_2 _3178_ (.A(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__o21ai_1 _3179_ (.A1(_2355_),
    .A2(_0695_),
    .B1(_0659_),
    .Y(_0696_));
 sky130_fd_sc_hd__nand2_1 _3180_ (.A(_2359_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__o21ai_1 _3181_ (.A1(_2356_),
    .A2(_2358_),
    .B1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__nand2_1 _3182_ (.A(_2361_),
    .B(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__o211a_1 _3183_ (.A1(_2361_),
    .A2(_0698_),
    .B1(_0688_),
    .C1(_0699_),
    .X(_0491_));
 sky130_fd_sc_hd__buf_1 _3184_ (.A(_0693_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_2 _3185_ (.A(_0679_),
    .X(_0700_));
 sky130_fd_sc_hd__clkbuf_2 _3186_ (.A(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__o211a_1 _3187_ (.A1(_2359_),
    .A2(_0696_),
    .B1(_0701_),
    .C1(_0697_),
    .X(_0490_));
 sky130_fd_sc_hd__buf_1 _3188_ (.A(_0693_),
    .X(_0139_));
 sky130_fd_sc_hd__or2_1 _3189_ (.A(_2349_),
    .B(_0695_),
    .X(_0702_));
 sky130_fd_sc_hd__o21ai_1 _3190_ (.A1(_2346_),
    .A2(_2347_),
    .B1(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__inv_2 _3191_ (.A(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__clkbuf_2 _3192_ (.A(_0680_),
    .X(_0705_));
 sky130_fd_sc_hd__buf_2 _3193_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__o221a_1 _3194_ (.A1(_2354_),
    .A2(_0704_),
    .B1(_2353_),
    .B2(_0703_),
    .C1(_0706_),
    .X(_0489_));
 sky130_fd_sc_hd__buf_1 _3195_ (.A(_0693_),
    .X(_0138_));
 sky130_fd_sc_hd__o211a_1 _3196_ (.A1(_2348_),
    .A2(_0694_),
    .B1(_0701_),
    .C1(_0702_),
    .X(_0488_));
 sky130_fd_sc_hd__buf_1 _3197_ (.A(_0693_),
    .X(_0137_));
 sky130_fd_sc_hd__o21ai_1 _3198_ (.A1(_0657_),
    .A2(_0511_),
    .B1(_0661_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand2_1 _3199_ (.A(_0500_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__o21ai_1 _3200_ (.A1(_2368_),
    .A2(_0499_),
    .B1(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _3201_ (.A(_2367_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o211a_1 _3202_ (.A1(_2367_),
    .A2(_0709_),
    .B1(_0701_),
    .C1(_0710_),
    .X(_0487_));
 sky130_fd_sc_hd__buf_1 _3203_ (.A(_2326_),
    .X(_0711_));
 sky130_fd_sc_hd__buf_1 _3204_ (.A(_0711_),
    .X(_0136_));
 sky130_fd_sc_hd__o211a_1 _3205_ (.A1(_0500_),
    .A2(_0707_),
    .B1(_0701_),
    .C1(_0708_),
    .X(_0486_));
 sky130_fd_sc_hd__buf_1 _3206_ (.A(_0711_),
    .X(_0135_));
 sky130_fd_sc_hd__or2_1 _3207_ (.A(_0657_),
    .B(_0510_),
    .X(_0712_));
 sky130_fd_sc_hd__o21ai_1 _3208_ (.A1(_0507_),
    .A2(_0508_),
    .B1(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__inv_2 _3209_ (.A(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__o221a_1 _3210_ (.A1(_0506_),
    .A2(_0714_),
    .B1(_0505_),
    .B2(_0713_),
    .C1(_0706_),
    .X(_0485_));
 sky130_fd_sc_hd__buf_1 _3211_ (.A(_0711_),
    .X(_0134_));
 sky130_fd_sc_hd__inv_2 _3212_ (.A(_0657_),
    .Y(_0715_));
 sky130_fd_sc_hd__o211a_1 _3213_ (.A1(_0715_),
    .A2(_0509_),
    .B1(_0701_),
    .C1(_0712_),
    .X(_0484_));
 sky130_fd_sc_hd__buf_1 _3214_ (.A(_0711_),
    .X(_0133_));
 sky130_fd_sc_hd__o21ai_1 _3215_ (.A1(_0642_),
    .A2(_0652_),
    .B1(_0542_),
    .Y(_0716_));
 sky130_fd_sc_hd__inv_2 _3216_ (.A(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__o21ai_1 _3217_ (.A1(_0528_),
    .A2(_0717_),
    .B1(_0545_),
    .Y(_0718_));
 sky130_fd_sc_hd__nand2_1 _3218_ (.A(_0655_),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__o21ai_1 _3219_ (.A1(_0516_),
    .A2(_0518_),
    .B1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__inv_2 _3220_ (.A(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__o221a_1 _3221_ (.A1(_0654_),
    .A2(_0721_),
    .B1(_0653_),
    .B2(_0720_),
    .C1(_0706_),
    .X(_0483_));
 sky130_fd_sc_hd__buf_1 _3222_ (.A(_0711_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_2 _3223_ (.A(_0700_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_1 _3224_ (.A1(_0655_),
    .A2(_0718_),
    .B1(_0722_),
    .C1(_0719_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_1 _3225_ (.A(_2326_),
    .X(_0723_));
 sky130_fd_sc_hd__buf_1 _3226_ (.A(_0723_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _3227_ (.A(_0527_),
    .B(_0717_),
    .X(_0724_));
 sky130_fd_sc_hd__o21ai_1 _3228_ (.A1(_0524_),
    .A2(_0525_),
    .B1(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__inv_2 _3229_ (.A(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__o221a_1 _3230_ (.A1(_0523_),
    .A2(_0726_),
    .B1(_0522_),
    .B2(_0725_),
    .C1(_0706_),
    .X(_0481_));
 sky130_fd_sc_hd__buf_1 _3231_ (.A(_0723_),
    .X(_0130_));
 sky130_fd_sc_hd__o211a_1 _3232_ (.A1(_0526_),
    .A2(_0716_),
    .B1(_0722_),
    .C1(_0724_),
    .X(_0480_));
 sky130_fd_sc_hd__buf_1 _3233_ (.A(_0723_),
    .X(_0129_));
 sky130_fd_sc_hd__o21ai_1 _3234_ (.A1(_0642_),
    .A2(_0651_),
    .B1(_0540_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _3235_ (.A(_0536_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__o21ai_1 _3236_ (.A1(_0533_),
    .A2(_0535_),
    .B1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__nand2_1 _3237_ (.A(_0532_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__o211a_1 _3238_ (.A1(_0532_),
    .A2(_0729_),
    .B1(_0722_),
    .C1(_0730_),
    .X(_0479_));
 sky130_fd_sc_hd__buf_1 _3239_ (.A(_0723_),
    .X(_0128_));
 sky130_fd_sc_hd__o211a_1 _3240_ (.A1(_0536_),
    .A2(_0727_),
    .B1(_0722_),
    .C1(_0728_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_1 _3241_ (.A(_0723_),
    .X(_0127_));
 sky130_fd_sc_hd__or2_1 _3242_ (.A(_0642_),
    .B(_0650_),
    .X(_0731_));
 sky130_fd_sc_hd__o21ai_1 _3243_ (.A1(_0647_),
    .A2(_0648_),
    .B1(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__inv_2 _3244_ (.A(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__o221a_1 _3245_ (.A1(_0646_),
    .A2(_0733_),
    .B1(_0645_),
    .B2(_0732_),
    .C1(_0706_),
    .X(_0477_));
 sky130_fd_sc_hd__buf_1 _3246_ (.A(net40),
    .X(_0734_));
 sky130_fd_sc_hd__buf_1 _3247_ (.A(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__buf_1 _3248_ (.A(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__buf_1 _3249_ (.A(_0736_),
    .X(_0126_));
 sky130_fd_sc_hd__inv_2 _3250_ (.A(_0642_),
    .Y(_0737_));
 sky130_fd_sc_hd__o211a_1 _3251_ (.A1(_0737_),
    .A2(_0649_),
    .B1(_0722_),
    .C1(_0731_),
    .X(_0476_));
 sky130_fd_sc_hd__buf_1 _3252_ (.A(_0736_),
    .X(_0125_));
 sky130_fd_sc_hd__o21ai_1 _3253_ (.A1(_0631_),
    .A2(_0585_),
    .B1(_0637_),
    .Y(_0738_));
 sky130_fd_sc_hd__inv_2 _3254_ (.A(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__o21ai_1 _3255_ (.A1(_0564_),
    .A2(_0739_),
    .B1(_0633_),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _3256_ (.A(_0553_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__o21ai_1 _3257_ (.A1(_0550_),
    .A2(_0552_),
    .B1(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__clkbuf_2 _3258_ (.A(_0700_),
    .X(_0743_));
 sky130_fd_sc_hd__nand2_1 _3259_ (.A(_0549_),
    .B(_0742_),
    .Y(_0744_));
 sky130_fd_sc_hd__o211a_1 _3260_ (.A1(_0549_),
    .A2(_0742_),
    .B1(_0743_),
    .C1(_0744_),
    .X(_0475_));
 sky130_fd_sc_hd__buf_1 _3261_ (.A(_0736_),
    .X(_0124_));
 sky130_fd_sc_hd__o211a_1 _3262_ (.A1(_0553_),
    .A2(_0740_),
    .B1(_0743_),
    .C1(_0741_),
    .X(_0474_));
 sky130_fd_sc_hd__buf_1 _3263_ (.A(_0736_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _3264_ (.A(_0563_),
    .B(_0739_),
    .X(_0745_));
 sky130_fd_sc_hd__o21ai_1 _3265_ (.A1(_0560_),
    .A2(_0561_),
    .B1(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__inv_2 _3266_ (.A(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__buf_2 _3267_ (.A(_0705_),
    .X(_0748_));
 sky130_fd_sc_hd__o221a_1 _3268_ (.A1(_0559_),
    .A2(_0747_),
    .B1(_0558_),
    .B2(_0746_),
    .C1(_0748_),
    .X(_0473_));
 sky130_fd_sc_hd__buf_1 _3269_ (.A(_0736_),
    .X(_0122_));
 sky130_fd_sc_hd__o211a_1 _3270_ (.A1(_0562_),
    .A2(_0738_),
    .B1(_0743_),
    .C1(_0745_),
    .X(_0472_));
 sky130_fd_sc_hd__buf_1 _3271_ (.A(_0735_),
    .X(_0749_));
 sky130_fd_sc_hd__buf_1 _3272_ (.A(_0749_),
    .X(_0121_));
 sky130_fd_sc_hd__o21ai_1 _3273_ (.A1(_0631_),
    .A2(_0584_),
    .B1(_0635_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2_1 _3274_ (.A(_0573_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__o21ai_1 _3275_ (.A1(_0570_),
    .A2(_0572_),
    .B1(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _3276_ (.A(_0569_),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__o211a_1 _3277_ (.A1(_0569_),
    .A2(_0752_),
    .B1(_0743_),
    .C1(_0753_),
    .X(_0471_));
 sky130_fd_sc_hd__buf_1 _3278_ (.A(_0749_),
    .X(_0120_));
 sky130_fd_sc_hd__o211a_1 _3279_ (.A1(_0573_),
    .A2(_0750_),
    .B1(_0743_),
    .C1(_0751_),
    .X(_0470_));
 sky130_fd_sc_hd__buf_1 _3280_ (.A(_0749_),
    .X(_0119_));
 sky130_fd_sc_hd__or2_1 _3281_ (.A(_0631_),
    .B(_0583_),
    .X(_0754_));
 sky130_fd_sc_hd__o21ai_1 _3282_ (.A1(_0580_),
    .A2(_0581_),
    .B1(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__inv_2 _3283_ (.A(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__o221a_1 _3284_ (.A1(_0579_),
    .A2(_0756_),
    .B1(_0578_),
    .B2(_0755_),
    .C1(_0748_),
    .X(_0469_));
 sky130_fd_sc_hd__buf_1 _3285_ (.A(_0749_),
    .X(_0118_));
 sky130_fd_sc_hd__inv_2 _3286_ (.A(_0631_),
    .Y(_0757_));
 sky130_fd_sc_hd__buf_2 _3287_ (.A(_0700_),
    .X(_0758_));
 sky130_fd_sc_hd__o211a_1 _3288_ (.A1(_0757_),
    .A2(_0582_),
    .B1(_0758_),
    .C1(_0754_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_1 _3289_ (.A(_0749_),
    .X(_0117_));
 sky130_fd_sc_hd__inv_2 _3290_ (.A(_0629_),
    .Y(_0759_));
 sky130_fd_sc_hd__a31o_1 _3291_ (.A1(_0605_),
    .A2(_0606_),
    .A3(_0759_),
    .B1(_0600_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_1 _3292_ (.A(_0592_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__o21ai_1 _3293_ (.A1(_0589_),
    .A2(_0591_),
    .B1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__inv_2 _3294_ (.A(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__o221a_1 _3295_ (.A1(_0588_),
    .A2(_0763_),
    .B1(_0587_),
    .B2(_0762_),
    .C1(_0748_),
    .X(_0467_));
 sky130_fd_sc_hd__buf_1 _3296_ (.A(_0735_),
    .X(_0764_));
 sky130_fd_sc_hd__buf_1 _3297_ (.A(_0764_),
    .X(_0116_));
 sky130_fd_sc_hd__o211a_1 _3298_ (.A1(_0592_),
    .A2(_0760_),
    .B1(_0758_),
    .C1(_0761_),
    .X(_0466_));
 sky130_fd_sc_hd__buf_1 _3299_ (.A(_0764_),
    .X(_0115_));
 sky130_fd_sc_hd__nand2_1 _3300_ (.A(_0759_),
    .B(_0606_),
    .Y(_0765_));
 sky130_fd_sc_hd__inv_2 _3301_ (.A(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__clkbuf_4 _3302_ (.A(_0681_),
    .X(_0767_));
 sky130_fd_sc_hd__o21ai_1 _3303_ (.A1(_0599_),
    .A2(_0766_),
    .B1(_0605_),
    .Y(_0768_));
 sky130_fd_sc_hd__o311a_1 _3304_ (.A1(_0599_),
    .A2(_0766_),
    .A3(_0605_),
    .B1(_0767_),
    .C1(_0768_),
    .X(_0465_));
 sky130_fd_sc_hd__buf_1 _3305_ (.A(_0764_),
    .X(_0114_));
 sky130_fd_sc_hd__o211a_1 _3306_ (.A1(_0759_),
    .A2(_0606_),
    .B1(_0758_),
    .C1(_0765_),
    .X(_0464_));
 sky130_fd_sc_hd__buf_1 _3307_ (.A(_0764_),
    .X(_0113_));
 sky130_fd_sc_hd__or2_1 _3308_ (.A(_0625_),
    .B(_0615_),
    .X(_0769_));
 sky130_fd_sc_hd__o21ai_1 _3309_ (.A1(_0611_),
    .A2(_0613_),
    .B1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__inv_2 _3310_ (.A(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__o221a_1 _3311_ (.A1(_0610_),
    .A2(_0771_),
    .B1(_0609_),
    .B2(_0770_),
    .C1(_0748_),
    .X(_0463_));
 sky130_fd_sc_hd__buf_1 _3312_ (.A(_0764_),
    .X(_0112_));
 sky130_fd_sc_hd__o211a_1 _3313_ (.A1(_0624_),
    .A2(_0614_),
    .B1(_0758_),
    .C1(_0769_),
    .X(_0462_));
 sky130_fd_sc_hd__buf_1 _3314_ (.A(_0735_),
    .X(_0772_));
 sky130_fd_sc_hd__buf_1 _3315_ (.A(_0772_),
    .X(_0111_));
 sky130_fd_sc_hd__o21a_1 _3316_ (.A1(_0619_),
    .A2(_0621_),
    .B1(_0622_),
    .X(_0773_));
 sky130_fd_sc_hd__clkbuf_2 _3317_ (.A(_0680_),
    .X(_0774_));
 sky130_fd_sc_hd__and3b_1 _3318_ (.A_N(_0773_),
    .B(_0623_),
    .C(_0774_),
    .X(_0461_));
 sky130_fd_sc_hd__buf_1 _3319_ (.A(_0772_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_2 _3320_ (.A(_0619_),
    .X(_0775_));
 sky130_fd_sc_hd__o221a_1 _3321_ (.A1(_0775_),
    .A2(_0621_),
    .B1(\acc1[0] ),
    .B2(\acc2[0] ),
    .C1(_0748_),
    .X(_0460_));
 sky130_fd_sc_hd__buf_1 _3322_ (.A(_0772_),
    .X(_0109_));
 sky130_fd_sc_hd__inv_1 _3323_ (.A(net17),
    .Y(_0776_));
 sky130_fd_sc_hd__or4_4 _3324_ (.A(_0619_),
    .B(_0776_),
    .C(_0616_),
    .D(_0611_),
    .X(_0777_));
 sky130_fd_sc_hd__or2_2 _3325_ (.A(_0626_),
    .B(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__or2_1 _3326_ (.A(_0597_),
    .B(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__or2_1 _3327_ (.A(_0594_),
    .B(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__or2_1 _3328_ (.A(_0589_),
    .B(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__or2_1 _3329_ (.A(_0602_),
    .B(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__or2_1 _3330_ (.A(_0580_),
    .B(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__or2_1 _3331_ (.A(_0575_),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__or2_1 _3332_ (.A(_0570_),
    .B(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__or2_1 _3333_ (.A(_0566_),
    .B(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__or2_1 _3334_ (.A(_0560_),
    .B(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__or2_1 _3335_ (.A(_0555_),
    .B(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__or2_1 _3336_ (.A(_0550_),
    .B(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__or2_1 _3337_ (.A(_0638_),
    .B(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__or2_1 _3338_ (.A(_0647_),
    .B(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__or2_1 _3339_ (.A(_0643_),
    .B(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__or2_1 _3340_ (.A(_0533_),
    .B(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__or2_1 _3341_ (.A(_0529_),
    .B(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__or2_1 _3342_ (.A(_0524_),
    .B(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__or2_1 _3343_ (.A(_0520_),
    .B(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__or2_2 _3344_ (.A(_0516_),
    .B(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__or2_2 _3345_ (.A(_0514_),
    .B(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__or2_1 _3346_ (.A(_0507_),
    .B(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__or2_1 _3347_ (.A(_0502_),
    .B(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__or2_1 _3348_ (.A(_2368_),
    .B(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__or2_1 _3349_ (.A(_2364_),
    .B(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__or2_1 _3350_ (.A(_2346_),
    .B(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__or2_1 _3351_ (.A(_2351_),
    .B(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__or2_1 _3352_ (.A(_2356_),
    .B(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__or2_1 _3353_ (.A(_0664_),
    .B(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__or2_1 _3354_ (.A(_2341_),
    .B(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__or2_1 _3355_ (.A(_0669_),
    .B(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__or2_2 _3356_ (.A(_2333_),
    .B(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__or2_4 _3357_ (.A(_0673_),
    .B(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__inv_2 _3358_ (.A(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__buf_2 _3359_ (.A(_0705_),
    .X(_0812_));
 sky130_fd_sc_hd__o221a_1 _3360_ (.A1(\acc1[36] ),
    .A2(_0811_),
    .B1(_2327_),
    .B2(_0810_),
    .C1(_0812_),
    .X(_0459_));
 sky130_fd_sc_hd__buf_1 _3361_ (.A(_0772_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_2 _3362_ (.A(net18),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_4 _3363_ (.A(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__a211oi_2 _3364_ (.A1(_0673_),
    .A2(net54),
    .B1(_0814_),
    .C1(_0811_),
    .Y(_0458_));
 sky130_fd_sc_hd__buf_1 _3365_ (.A(_0772_),
    .X(_0107_));
 sky130_fd_sc_hd__inv_2 _3366_ (.A(net94),
    .Y(_0815_));
 sky130_fd_sc_hd__o211a_1 _3367_ (.A1(\acc1[34] ),
    .A2(_0815_),
    .B1(_0758_),
    .C1(net53),
    .X(_0457_));
 sky130_fd_sc_hd__buf_1 _3368_ (.A(_0735_),
    .X(_0816_));
 sky130_fd_sc_hd__buf_1 _3369_ (.A(_0816_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_2 _3370_ (.A(net18),
    .X(_0817_));
 sky130_fd_sc_hd__buf_2 _3371_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__a211oi_1 _3372_ (.A1(_0669_),
    .A2(net69),
    .B1(_0818_),
    .C1(_0815_),
    .Y(_0456_));
 sky130_fd_sc_hd__buf_1 _3373_ (.A(_0816_),
    .X(_0105_));
 sky130_fd_sc_hd__inv_2 _3374_ (.A(net81),
    .Y(_0819_));
 sky130_fd_sc_hd__buf_2 _3375_ (.A(_0700_),
    .X(_0820_));
 sky130_fd_sc_hd__o211a_1 _3376_ (.A1(\acc1[32] ),
    .A2(_0819_),
    .B1(_0820_),
    .C1(net69),
    .X(_0455_));
 sky130_fd_sc_hd__buf_1 _3377_ (.A(_0816_),
    .X(_0104_));
 sky130_fd_sc_hd__a211oi_1 _3378_ (.A1(_0664_),
    .A2(net60),
    .B1(_0818_),
    .C1(_0819_),
    .Y(_0454_));
 sky130_fd_sc_hd__buf_1 _3379_ (.A(_0816_),
    .X(_0103_));
 sky130_fd_sc_hd__inv_2 _3380_ (.A(net90),
    .Y(_0821_));
 sky130_fd_sc_hd__o211a_1 _3381_ (.A1(\acc1[30] ),
    .A2(_0821_),
    .B1(_0820_),
    .C1(net59),
    .X(_0453_));
 sky130_fd_sc_hd__buf_1 _3382_ (.A(_0816_),
    .X(_0102_));
 sky130_fd_sc_hd__a211oi_1 _3383_ (.A1(_2351_),
    .A2(net49),
    .B1(_0818_),
    .C1(_0821_),
    .Y(_0452_));
 sky130_fd_sc_hd__buf_1 _3384_ (.A(_0734_),
    .X(_0822_));
 sky130_fd_sc_hd__buf_1 _3385_ (.A(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__buf_1 _3386_ (.A(_0823_),
    .X(_0101_));
 sky130_fd_sc_hd__clkinvlp_2 _3387_ (.A(net89),
    .Y(_0824_));
 sky130_fd_sc_hd__o211a_1 _3388_ (.A1(\acc1[28] ),
    .A2(_0824_),
    .B1(_0820_),
    .C1(net48),
    .X(_0451_));
 sky130_fd_sc_hd__buf_1 _3389_ (.A(_0823_),
    .X(_0100_));
 sky130_fd_sc_hd__a211oi_1 _3390_ (.A1(_2364_),
    .A2(net56),
    .B1(_0818_),
    .C1(_0824_),
    .Y(_0450_));
 sky130_fd_sc_hd__buf_1 _3391_ (.A(_0823_),
    .X(_0099_));
 sky130_fd_sc_hd__clkinvlp_2 _3392_ (.A(net78),
    .Y(_0825_));
 sky130_fd_sc_hd__o211a_1 _3393_ (.A1(\acc1[26] ),
    .A2(_0825_),
    .B1(_0820_),
    .C1(net55),
    .X(_0449_));
 sky130_fd_sc_hd__buf_1 _3394_ (.A(_0823_),
    .X(_0098_));
 sky130_fd_sc_hd__a211oi_1 _3395_ (.A1(_0502_),
    .A2(net80),
    .B1(_0818_),
    .C1(_0825_),
    .Y(_0448_));
 sky130_fd_sc_hd__buf_1 _3396_ (.A(_0823_),
    .X(_0097_));
 sky130_fd_sc_hd__inv_2 _3397_ (.A(net50),
    .Y(_0826_));
 sky130_fd_sc_hd__o211a_1 _3398_ (.A1(\acc1[24] ),
    .A2(_0826_),
    .B1(_0820_),
    .C1(net79),
    .X(_0447_));
 sky130_fd_sc_hd__buf_1 _3399_ (.A(_0822_),
    .X(_0827_));
 sky130_fd_sc_hd__buf_1 _3400_ (.A(_0827_),
    .X(_0096_));
 sky130_fd_sc_hd__buf_2 _3401_ (.A(_0817_),
    .X(_0828_));
 sky130_fd_sc_hd__a211oi_2 _3402_ (.A1(_0514_),
    .A2(net64),
    .B1(_0828_),
    .C1(_0826_),
    .Y(_0446_));
 sky130_fd_sc_hd__buf_1 _3403_ (.A(_0827_),
    .X(_0095_));
 sky130_fd_sc_hd__inv_2 _3404_ (.A(net91),
    .Y(_0829_));
 sky130_fd_sc_hd__clkbuf_4 _3405_ (.A(_0679_),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_2 _3406_ (.A(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__o211a_1 _3407_ (.A1(\acc1[22] ),
    .A2(_0829_),
    .B1(_0831_),
    .C1(net63),
    .X(_0445_));
 sky130_fd_sc_hd__buf_1 _3408_ (.A(_0827_),
    .X(_0094_));
 sky130_fd_sc_hd__a211oi_1 _3409_ (.A1(_0520_),
    .A2(net62),
    .B1(_0828_),
    .C1(_0829_),
    .Y(_0444_));
 sky130_fd_sc_hd__buf_1 _3410_ (.A(_0827_),
    .X(_0093_));
 sky130_fd_sc_hd__inv_2 _3411_ (.A(net93),
    .Y(_0832_));
 sky130_fd_sc_hd__o211a_1 _3412_ (.A1(\acc1[20] ),
    .A2(_0832_),
    .B1(_0831_),
    .C1(net61),
    .X(_0443_));
 sky130_fd_sc_hd__buf_1 _3413_ (.A(_0827_),
    .X(_0092_));
 sky130_fd_sc_hd__a211oi_1 _3414_ (.A1(_0529_),
    .A2(net58),
    .B1(_0828_),
    .C1(_0832_),
    .Y(_0442_));
 sky130_fd_sc_hd__buf_1 _3415_ (.A(_0822_),
    .X(_0833_));
 sky130_fd_sc_hd__buf_1 _3416_ (.A(_0833_),
    .X(_0091_));
 sky130_fd_sc_hd__clkinvlp_2 _3417_ (.A(net83),
    .Y(_0834_));
 sky130_fd_sc_hd__o211a_1 _3418_ (.A1(\acc1[18] ),
    .A2(_0834_),
    .B1(_0831_),
    .C1(net57),
    .X(_0441_));
 sky130_fd_sc_hd__buf_1 _3419_ (.A(_0833_),
    .X(_0090_));
 sky130_fd_sc_hd__a211oi_1 _3420_ (.A1(_0643_),
    .A2(net71),
    .B1(_0828_),
    .C1(_0834_),
    .Y(_0440_));
 sky130_fd_sc_hd__buf_1 _3421_ (.A(_0833_),
    .X(_0089_));
 sky130_fd_sc_hd__clkinvlp_2 _3422_ (.A(net77),
    .Y(_0835_));
 sky130_fd_sc_hd__o211a_1 _3423_ (.A1(\acc1[16] ),
    .A2(_0835_),
    .B1(_0831_),
    .C1(net70),
    .X(_0439_));
 sky130_fd_sc_hd__buf_1 _3424_ (.A(_0833_),
    .X(_0088_));
 sky130_fd_sc_hd__a211oi_1 _3425_ (.A1(_0638_),
    .A2(net88),
    .B1(_0828_),
    .C1(_0835_),
    .Y(_0438_));
 sky130_fd_sc_hd__buf_1 _3426_ (.A(_0833_),
    .X(_0087_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(net74),
    .Y(_0836_));
 sky130_fd_sc_hd__o211a_1 _3428_ (.A1(\acc1[14] ),
    .A2(_0836_),
    .B1(_0831_),
    .C1(net87),
    .X(_0437_));
 sky130_fd_sc_hd__buf_1 _3429_ (.A(_0822_),
    .X(_0837_));
 sky130_fd_sc_hd__buf_1 _3430_ (.A(_0837_),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_2 _3431_ (.A(_0813_),
    .X(_0838_));
 sky130_fd_sc_hd__a211oi_1 _3432_ (.A1(_0555_),
    .A2(net76),
    .B1(_0838_),
    .C1(_0836_),
    .Y(_0436_));
 sky130_fd_sc_hd__buf_1 _3433_ (.A(_0837_),
    .X(_0085_));
 sky130_fd_sc_hd__inv_2 _3434_ (.A(net92),
    .Y(_0839_));
 sky130_fd_sc_hd__clkbuf_2 _3435_ (.A(_0830_),
    .X(_0840_));
 sky130_fd_sc_hd__o211a_1 _3436_ (.A1(\acc1[12] ),
    .A2(_0839_),
    .B1(_0840_),
    .C1(net75),
    .X(_0435_));
 sky130_fd_sc_hd__buf_1 _3437_ (.A(_0837_),
    .X(_0084_));
 sky130_fd_sc_hd__a211oi_1 _3438_ (.A1(_0566_),
    .A2(net68),
    .B1(_0838_),
    .C1(_0839_),
    .Y(_0434_));
 sky130_fd_sc_hd__buf_1 _3439_ (.A(_0837_),
    .X(_0083_));
 sky130_fd_sc_hd__inv_2 _3440_ (.A(net86),
    .Y(_0841_));
 sky130_fd_sc_hd__o211a_1 _3441_ (.A1(\acc1[10] ),
    .A2(_0841_),
    .B1(_0840_),
    .C1(net67),
    .X(_0433_));
 sky130_fd_sc_hd__buf_1 _3442_ (.A(_0837_),
    .X(_0082_));
 sky130_fd_sc_hd__a211oi_1 _3443_ (.A1(_0575_),
    .A2(net73),
    .B1(_0838_),
    .C1(_0841_),
    .Y(_0432_));
 sky130_fd_sc_hd__buf_1 _3444_ (.A(_0822_),
    .X(_0842_));
 sky130_fd_sc_hd__buf_1 _3445_ (.A(_0842_),
    .X(_0081_));
 sky130_fd_sc_hd__inv_2 _3446_ (.A(net84),
    .Y(_0843_));
 sky130_fd_sc_hd__o211a_1 _3447_ (.A1(\acc1[8] ),
    .A2(_0843_),
    .B1(_0840_),
    .C1(net72),
    .X(_0431_));
 sky130_fd_sc_hd__buf_1 _3448_ (.A(_0842_),
    .X(_0080_));
 sky130_fd_sc_hd__a211oi_1 _3449_ (.A1(_0602_),
    .A2(net66),
    .B1(_0838_),
    .C1(_0843_),
    .Y(_0430_));
 sky130_fd_sc_hd__buf_1 _3450_ (.A(_0842_),
    .X(_0079_));
 sky130_fd_sc_hd__inv_2 _3451_ (.A(net82),
    .Y(_0844_));
 sky130_fd_sc_hd__o211a_1 _3452_ (.A1(\acc1[6] ),
    .A2(_0844_),
    .B1(_0840_),
    .C1(net65),
    .X(_0429_));
 sky130_fd_sc_hd__buf_1 _3453_ (.A(_0842_),
    .X(_0078_));
 sky130_fd_sc_hd__a211oi_2 _3454_ (.A1(_0594_),
    .A2(net51),
    .B1(_0838_),
    .C1(_0844_),
    .Y(_0428_));
 sky130_fd_sc_hd__buf_1 _3455_ (.A(_0842_),
    .X(_0077_));
 sky130_fd_sc_hd__inv_2 _3456_ (.A(net43),
    .Y(_0845_));
 sky130_fd_sc_hd__o211a_1 _3457_ (.A1(\acc1[4] ),
    .A2(_0845_),
    .B1(_0840_),
    .C1(net52),
    .X(_0427_));
 sky130_fd_sc_hd__buf_1 _3458_ (.A(net39),
    .X(_0846_));
 sky130_fd_sc_hd__buf_1 _3459_ (.A(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_1 _3460_ (.A(_0847_),
    .X(_0076_));
 sky130_fd_sc_hd__inv_2 _3461_ (.A(_0777_),
    .Y(_0848_));
 sky130_fd_sc_hd__buf_2 _3462_ (.A(_0830_),
    .X(_0849_));
 sky130_fd_sc_hd__o211a_1 _3463_ (.A1(\acc1[3] ),
    .A2(_0848_),
    .B1(_0849_),
    .C1(net42),
    .X(_0426_));
 sky130_fd_sc_hd__buf_1 _3464_ (.A(_0847_),
    .X(_0075_));
 sky130_fd_sc_hd__o31a_1 _3465_ (.A1(_0775_),
    .A2(net47),
    .A3(_0617_),
    .B1(_0611_),
    .X(_0850_));
 sky130_fd_sc_hd__nor3_1 _3466_ (.A(_0814_),
    .B(_0848_),
    .C(_0850_),
    .Y(_0425_));
 sky130_fd_sc_hd__buf_1 _3467_ (.A(_0847_),
    .X(_0074_));
 sky130_fd_sc_hd__o21ai_1 _3468_ (.A1(_0775_),
    .A2(net46),
    .B1(_0617_),
    .Y(_0851_));
 sky130_fd_sc_hd__o311a_1 _3469_ (.A1(_0775_),
    .A2(net45),
    .A3(_0617_),
    .B1(_0767_),
    .C1(_0851_),
    .X(_0424_));
 sky130_fd_sc_hd__buf_1 _3470_ (.A(_0847_),
    .X(_0073_));
 sky130_fd_sc_hd__o221a_1 _3471_ (.A1(_0775_),
    .A2(net44),
    .B1(\acc1[0] ),
    .B2(net85),
    .C1(_0812_),
    .X(_0423_));
 sky130_fd_sc_hd__inv_2 _3472_ (.A(\word_count[12] ),
    .Y(_0852_));
 sky130_fd_sc_hd__inv_2 _3473_ (.A(\word_count[10] ),
    .Y(_0853_));
 sky130_fd_sc_hd__and3_1 _3474_ (.A(\word_count[0] ),
    .B(\word_count[1] ),
    .C(\word_count[2] ),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _3475_ (.A(\word_count[3] ),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__inv_2 _3476_ (.A(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand2_1 _3477_ (.A(\word_count[4] ),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__or2_1 _3478_ (.A(_2294_),
    .B(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__or2_2 _3479_ (.A(_2285_),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__nor2_2 _3480_ (.A(_2291_),
    .B(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__nand2_1 _3481_ (.A(_2272_),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__inv_2 _3482_ (.A(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__nand2_1 _3483_ (.A(_2270_),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__or2_1 _3484_ (.A(_0853_),
    .B(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__or2_1 _3485_ (.A(_2278_),
    .B(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__or2_1 _3486_ (.A(_0852_),
    .B(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__or2_1 _3487_ (.A(_2276_),
    .B(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__or2_1 _3488_ (.A(_2244_),
    .B(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__inv_2 _3489_ (.A(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__inv_2 _3490_ (.A(net7),
    .Y(_0870_));
 sky130_fd_sc_hd__clkbuf_2 _3491_ (.A(net1),
    .X(_0871_));
 sky130_fd_sc_hd__buf_1 _3492_ (.A(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__clkbuf_2 _3493_ (.A(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__nor2_1 _3494_ (.A(_0873_),
    .B(_2256_),
    .Y(_0874_));
 sky130_fd_sc_hd__o22a_1 _3495_ (.A1(_0870_),
    .A2(_0874_),
    .B1(_0873_),
    .B2(_2259_),
    .X(_0875_));
 sky130_fd_sc_hd__inv_2 _3496_ (.A(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__o22a_1 _3497_ (.A1(_2281_),
    .A2(_0875_),
    .B1(\word_count[15] ),
    .B2(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__or2_1 _3498_ (.A(_0873_),
    .B(_2255_),
    .X(_0878_));
 sky130_fd_sc_hd__a21oi_2 _3499_ (.A1(net6),
    .A2(_0878_),
    .B1(_0874_),
    .Y(_0879_));
 sky130_fd_sc_hd__inv_2 _3500_ (.A(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__inv_2 _3501_ (.A(net16),
    .Y(_0881_));
 sky130_fd_sc_hd__nor2_1 _3502_ (.A(_0872_),
    .B(_2251_),
    .Y(_0882_));
 sky130_fd_sc_hd__or2_1 _3503_ (.A(_0872_),
    .B(_2252_),
    .X(_0883_));
 sky130_fd_sc_hd__o21a_1 _3504_ (.A1(_0881_),
    .A2(_0882_),
    .B1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__a2bb2o_1 _3505_ (.A1_N(_2270_),
    .A2_N(_0884_),
    .B1(\word_count[9] ),
    .B2(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__inv_2 _3506_ (.A(net4),
    .Y(_0886_));
 sky130_fd_sc_hd__nor2_1 _3507_ (.A(_0872_),
    .B(_2258_),
    .Y(_0887_));
 sky130_fd_sc_hd__or2_1 _3508_ (.A(_0872_),
    .B(_2254_),
    .X(_0888_));
 sky130_fd_sc_hd__o21a_1 _3509_ (.A1(_0886_),
    .A2(_0887_),
    .B1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__a2bb2o_1 _3510_ (.A1_N(\word_count[12] ),
    .A2_N(_0889_),
    .B1(\word_count[12] ),
    .B2(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__inv_2 _3511_ (.A(_0871_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_1 _3512_ (.A(_0891_),
    .B(_2267_),
    .Y(_0892_));
 sky130_fd_sc_hd__inv_2 _3513_ (.A(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__o22a_1 _3514_ (.A1(_2265_),
    .A2(_0892_),
    .B1(net3),
    .B2(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__or2_2 _3515_ (.A(_0871_),
    .B(_2247_),
    .X(_0895_));
 sky130_fd_sc_hd__or2_1 _3516_ (.A(net12),
    .B(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__or2_2 _3517_ (.A(_2292_),
    .B(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__or2_1 _3518_ (.A(_0871_),
    .B(_2250_),
    .X(_0898_));
 sky130_fd_sc_hd__a21bo_1 _3519_ (.A1(net14),
    .A2(_0897_),
    .B1_N(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__o2bb2a_1 _3520_ (.A1_N(\word_count[7] ),
    .A2_N(_0899_),
    .B1(\word_count[7] ),
    .B2(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__or2_1 _3521_ (.A(net1),
    .B(net8),
    .X(_0901_));
 sky130_fd_sc_hd__or2_1 _3522_ (.A(net9),
    .B(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__nor2_1 _3523_ (.A(net10),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__a21oi_1 _3524_ (.A1(net10),
    .A2(_0902_),
    .B1(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor2_1 _3525_ (.A(_2307_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__o22a_1 _3526_ (.A1(_2300_),
    .A2(_0871_),
    .B1(\word_count[0] ),
    .B2(_0891_),
    .X(_0906_));
 sky130_fd_sc_hd__o21ai_1 _3527_ (.A1(_2300_),
    .A2(net8),
    .B1(_2304_),
    .Y(_0907_));
 sky130_fd_sc_hd__o2bb2a_1 _3528_ (.A1_N(\word_count[1] ),
    .A2_N(_0907_),
    .B1(\word_count[1] ),
    .B2(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__a21bo_1 _3529_ (.A1(net9),
    .A2(_0901_),
    .B1_N(_0902_),
    .X(_0909_));
 sky130_fd_sc_hd__a2bb2o_1 _3530_ (.A1_N(_2296_),
    .A2_N(_0909_),
    .B1(_2296_),
    .B2(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__or3_1 _3531_ (.A(_0906_),
    .B(_0908_),
    .C(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__inv_2 _3532_ (.A(net11),
    .Y(_0912_));
 sky130_fd_sc_hd__o21a_1 _3533_ (.A1(_0912_),
    .A2(_0903_),
    .B1(_0895_),
    .X(_0913_));
 sky130_fd_sc_hd__a2bb2o_1 _3534_ (.A1_N(_2311_),
    .A2_N(_0913_),
    .B1(_2311_),
    .B2(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__a2111o_1 _3535_ (.A1(_2307_),
    .A2(_0904_),
    .B1(_0905_),
    .C1(_0911_),
    .D1(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a21boi_1 _3536_ (.A1(net12),
    .A2(_0895_),
    .B1_N(_0896_),
    .Y(_0916_));
 sky130_fd_sc_hd__a2bb2o_1 _3537_ (.A1_N(\word_count[5] ),
    .A2_N(_0916_),
    .B1(\word_count[5] ),
    .B2(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__a21bo_1 _3538_ (.A1(_2292_),
    .A2(_0896_),
    .B1_N(_0897_),
    .X(_0918_));
 sky130_fd_sc_hd__a2bb2o_1 _3539_ (.A1_N(_2285_),
    .A2_N(_0918_),
    .B1(_2285_),
    .B2(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__a21oi_1 _3540_ (.A1(net15),
    .A2(_0898_),
    .B1(_0882_),
    .Y(_0920_));
 sky130_fd_sc_hd__a2bb2o_1 _3541_ (.A1_N(_2272_),
    .A2_N(_0920_),
    .B1(\word_count[8] ),
    .B2(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__or4_4 _3542_ (.A(_0915_),
    .B(_0917_),
    .C(_0919_),
    .D(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__a211o_1 _3543_ (.A1(_2278_),
    .A2(_0894_),
    .B1(_0900_),
    .C1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__or3_1 _3544_ (.A(_0885_),
    .B(_0890_),
    .C(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__a221o_1 _3545_ (.A1(\word_count[14] ),
    .A2(_0879_),
    .B1(_2244_),
    .B2(_0880_),
    .C1(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__a21boi_1 _3546_ (.A1(net5),
    .A2(_0888_),
    .B1_N(_0878_),
    .Y(_0926_));
 sky130_fd_sc_hd__a21oi_1 _3547_ (.A1(_2266_),
    .A2(_0883_),
    .B1(_0893_),
    .Y(_0927_));
 sky130_fd_sc_hd__a2bb2o_1 _3548_ (.A1_N(\word_count[10] ),
    .A2_N(_0927_),
    .B1(\word_count[10] ),
    .B2(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__a21oi_1 _3549_ (.A1(\word_count[13] ),
    .A2(_0926_),
    .B1(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__o221a_1 _3550_ (.A1(\word_count[13] ),
    .A2(_0926_),
    .B1(_2278_),
    .B2(_0894_),
    .C1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__or3b_2 _3551_ (.A(_0877_),
    .B(_0925_),
    .C_N(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__o21ba_2 _3552_ (.A1(_2263_),
    .A2(_2322_),
    .B1_N(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__inv_2 _3553_ (.A(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__clkbuf_2 _3554_ (.A(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__o221a_1 _3555_ (.A1(\word_count[15] ),
    .A2(_0869_),
    .B1(_2281_),
    .B2(_0868_),
    .C1(_0934_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_2 _3556_ (.A(_0932_),
    .X(_0030_));
 sky130_fd_sc_hd__a211oi_1 _3557_ (.A1(_2244_),
    .A2(_0867_),
    .B1(_0869_),
    .C1(_0030_),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_2 _3558_ (.A(_0866_),
    .Y(_0935_));
 sky130_fd_sc_hd__clkbuf_2 _3559_ (.A(_0933_),
    .X(_0936_));
 sky130_fd_sc_hd__o211a_1 _3560_ (.A1(\word_count[13] ),
    .A2(_0935_),
    .B1(_0867_),
    .C1(_0936_),
    .X(_0420_));
 sky130_fd_sc_hd__a211oi_1 _3561_ (.A1(_0852_),
    .A2(_0865_),
    .B1(_0935_),
    .C1(_0030_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_2 _3562_ (.A(_0864_),
    .Y(_0937_));
 sky130_fd_sc_hd__o211a_1 _3563_ (.A1(\word_count[11] ),
    .A2(_0937_),
    .B1(_0865_),
    .C1(_0936_),
    .X(_0418_));
 sky130_fd_sc_hd__a211oi_1 _3564_ (.A1(_0853_),
    .A2(_0863_),
    .B1(_0937_),
    .C1(_0932_),
    .Y(_0417_));
 sky130_fd_sc_hd__o211a_1 _3565_ (.A1(_2270_),
    .A2(_0862_),
    .B1(_0863_),
    .C1(_0936_),
    .X(_0416_));
 sky130_fd_sc_hd__o211a_1 _3566_ (.A1(_2272_),
    .A2(_0860_),
    .B1(_0861_),
    .C1(_0936_),
    .X(_0415_));
 sky130_fd_sc_hd__a211oi_2 _3567_ (.A1(_2291_),
    .A2(_0859_),
    .B1(_0860_),
    .C1(_0932_),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_2 _3568_ (.A(_0858_),
    .Y(_0938_));
 sky130_fd_sc_hd__o211a_1 _3569_ (.A1(\word_count[6] ),
    .A2(_0938_),
    .B1(_0859_),
    .C1(_0936_),
    .X(_0413_));
 sky130_fd_sc_hd__a211oi_2 _3570_ (.A1(_2294_),
    .A2(_0857_),
    .B1(_0938_),
    .C1(_0932_),
    .Y(_0412_));
 sky130_fd_sc_hd__o211a_1 _3571_ (.A1(_2311_),
    .A2(_0856_),
    .B1(_0857_),
    .C1(_0934_),
    .X(_0411_));
 sky130_fd_sc_hd__o211a_1 _3572_ (.A1(_2307_),
    .A2(_0854_),
    .B1(_0855_),
    .C1(_0934_),
    .X(_0410_));
 sky130_fd_sc_hd__o21a_1 _3573_ (.A1(_2300_),
    .A2(_2301_),
    .B1(_2296_),
    .X(_0939_));
 sky130_fd_sc_hd__nor3_1 _3574_ (.A(_0854_),
    .B(_0939_),
    .C(_0030_),
    .Y(_0409_));
 sky130_fd_sc_hd__o221a_1 _3575_ (.A1(_2300_),
    .A2(_2301_),
    .B1(\word_count[0] ),
    .B2(\word_count[1] ),
    .C1(_0934_),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_1 _3576_ (.A(\word_count[0] ),
    .B(_0030_),
    .Y(_0407_));
 sky130_fd_sc_hd__and2_1 _3577_ (.A(_0682_),
    .B(\diff2[36] ),
    .X(_0406_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3578_ (.A(_2324_),
    .X(_0940_));
 sky130_fd_sc_hd__inv_2 _3579_ (.A(\diff2[35] ),
    .Y(_0941_));
 sky130_fd_sc_hd__nor2_1 _3580_ (.A(_0940_),
    .B(_0941_),
    .Y(_0405_));
 sky130_fd_sc_hd__inv_2 _3581_ (.A(\diff2[34] ),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_1 _3582_ (.A(_0940_),
    .B(_0942_),
    .Y(_0404_));
 sky130_fd_sc_hd__inv_2 _3583_ (.A(\diff2[33] ),
    .Y(_0943_));
 sky130_fd_sc_hd__nor2_1 _3584_ (.A(_0940_),
    .B(_0943_),
    .Y(_0403_));
 sky130_fd_sc_hd__inv_2 _3585_ (.A(\diff2[32] ),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_1 _3586_ (.A(_0940_),
    .B(_0944_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _3587_ (.A(\diff2[31] ),
    .Y(_0945_));
 sky130_fd_sc_hd__nor2_1 _3588_ (.A(_0940_),
    .B(_0945_),
    .Y(_0401_));
 sky130_fd_sc_hd__clkbuf_2 _3589_ (.A(_2324_),
    .X(_0946_));
 sky130_fd_sc_hd__inv_2 _3590_ (.A(\diff2[30] ),
    .Y(_0947_));
 sky130_fd_sc_hd__nor2_1 _3591_ (.A(_0946_),
    .B(_0947_),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_2 _3592_ (.A(\diff2[29] ),
    .Y(_0948_));
 sky130_fd_sc_hd__nor2_1 _3593_ (.A(_0946_),
    .B(_0948_),
    .Y(_0399_));
 sky130_fd_sc_hd__inv_2 _3594_ (.A(\diff2[28] ),
    .Y(_0949_));
 sky130_fd_sc_hd__nor2_1 _3595_ (.A(_0946_),
    .B(_0949_),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _3596_ (.A(\diff2[27] ),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_1 _3597_ (.A(_0946_),
    .B(_0950_),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_2 _3598_ (.A(\diff2[26] ),
    .Y(_0951_));
 sky130_fd_sc_hd__nor2_1 _3599_ (.A(_0946_),
    .B(_0951_),
    .Y(_0396_));
 sky130_fd_sc_hd__clkbuf_2 _3600_ (.A(_2324_),
    .X(_0952_));
 sky130_fd_sc_hd__inv_2 _3601_ (.A(\diff2[25] ),
    .Y(_0953_));
 sky130_fd_sc_hd__nor2_1 _3602_ (.A(_0952_),
    .B(_0953_),
    .Y(_0395_));
 sky130_fd_sc_hd__inv_2 _3603_ (.A(\diff2[24] ),
    .Y(_0954_));
 sky130_fd_sc_hd__nor2_1 _3604_ (.A(_0952_),
    .B(_0954_),
    .Y(_0394_));
 sky130_fd_sc_hd__inv_2 _3605_ (.A(\diff2[23] ),
    .Y(_0955_));
 sky130_fd_sc_hd__nor2_1 _3606_ (.A(_0952_),
    .B(_0955_),
    .Y(_0393_));
 sky130_fd_sc_hd__inv_2 _3607_ (.A(\diff2[22] ),
    .Y(_0956_));
 sky130_fd_sc_hd__buf_1 _3608_ (.A(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__nor2_1 _3609_ (.A(_0952_),
    .B(_0957_),
    .Y(_0392_));
 sky130_fd_sc_hd__inv_2 _3610_ (.A(\diff2[21] ),
    .Y(_0958_));
 sky130_fd_sc_hd__nor2_1 _3611_ (.A(_0952_),
    .B(_0958_),
    .Y(_0391_));
 sky130_fd_sc_hd__buf_1 _3612_ (.A(_2324_),
    .X(_0959_));
 sky130_fd_sc_hd__inv_2 _3613_ (.A(\diff2[20] ),
    .Y(_0960_));
 sky130_fd_sc_hd__nor2_1 _3614_ (.A(_0959_),
    .B(_0960_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _3615_ (.A(\diff2[19] ),
    .Y(_0961_));
 sky130_fd_sc_hd__nor2_1 _3616_ (.A(_0959_),
    .B(_0961_),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_2 _3617_ (.A(\diff2[18] ),
    .Y(_0962_));
 sky130_fd_sc_hd__nor2_1 _3618_ (.A(_0959_),
    .B(_0962_),
    .Y(_0388_));
 sky130_fd_sc_hd__inv_2 _3619_ (.A(\diff2[17] ),
    .Y(_0963_));
 sky130_fd_sc_hd__nor2_1 _3620_ (.A(_0959_),
    .B(_0963_),
    .Y(_0387_));
 sky130_fd_sc_hd__inv_2 _3621_ (.A(\diff2[16] ),
    .Y(_0964_));
 sky130_fd_sc_hd__nor2_1 _3622_ (.A(_0959_),
    .B(_0964_),
    .Y(_0386_));
 sky130_fd_sc_hd__buf_2 _3623_ (.A(_0813_),
    .X(_0965_));
 sky130_fd_sc_hd__clkbuf_2 _3624_ (.A(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__inv_2 _3625_ (.A(\diff2[15] ),
    .Y(_0967_));
 sky130_fd_sc_hd__nor2_1 _3626_ (.A(_0966_),
    .B(_0967_),
    .Y(_0385_));
 sky130_fd_sc_hd__inv_2 _3627_ (.A(\diff2[14] ),
    .Y(_0968_));
 sky130_fd_sc_hd__nor2_1 _3628_ (.A(_0966_),
    .B(_0968_),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_2 _3629_ (.A(\diff2[13] ),
    .Y(_0969_));
 sky130_fd_sc_hd__nor2_1 _3630_ (.A(_0966_),
    .B(_0969_),
    .Y(_0383_));
 sky130_fd_sc_hd__inv_2 _3631_ (.A(\diff2[12] ),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_1 _3632_ (.A(_0966_),
    .B(_0970_),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_2 _3633_ (.A(\diff2[11] ),
    .Y(_0971_));
 sky130_fd_sc_hd__nor2_1 _3634_ (.A(_0966_),
    .B(_0971_),
    .Y(_0381_));
 sky130_fd_sc_hd__clkbuf_2 _3635_ (.A(_0965_),
    .X(_0972_));
 sky130_fd_sc_hd__inv_2 _3636_ (.A(\diff2[10] ),
    .Y(_0973_));
 sky130_fd_sc_hd__nor2_1 _3637_ (.A(_0972_),
    .B(_0973_),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _3638_ (.A(\diff2[9] ),
    .Y(_0974_));
 sky130_fd_sc_hd__nor2_1 _3639_ (.A(_0972_),
    .B(_0974_),
    .Y(_0379_));
 sky130_fd_sc_hd__inv_2 _3640_ (.A(\diff2[8] ),
    .Y(_0975_));
 sky130_fd_sc_hd__nor2_1 _3641_ (.A(_0972_),
    .B(_0975_),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(\diff2[7] ),
    .Y(_0976_));
 sky130_fd_sc_hd__nor2_1 _3643_ (.A(_0972_),
    .B(_0976_),
    .Y(_0377_));
 sky130_fd_sc_hd__inv_2 _3644_ (.A(\diff2[6] ),
    .Y(_0977_));
 sky130_fd_sc_hd__nor2_1 _3645_ (.A(_0972_),
    .B(_0977_),
    .Y(_0376_));
 sky130_fd_sc_hd__clkbuf_2 _3646_ (.A(_0965_),
    .X(_0978_));
 sky130_fd_sc_hd__inv_2 _3647_ (.A(\diff2[5] ),
    .Y(_0979_));
 sky130_fd_sc_hd__nor2_1 _3648_ (.A(_0978_),
    .B(_0979_),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_2 _3649_ (.A(\diff2[4] ),
    .Y(_0980_));
 sky130_fd_sc_hd__nor2_1 _3650_ (.A(_0978_),
    .B(_0980_),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(\diff2[3] ),
    .Y(_0981_));
 sky130_fd_sc_hd__nor2_1 _3652_ (.A(_0978_),
    .B(_0981_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _3653_ (.A(\diff2[2] ),
    .Y(_0982_));
 sky130_fd_sc_hd__nor2_1 _3654_ (.A(_0978_),
    .B(_0982_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _3655_ (.A(\diff2[1] ),
    .Y(_0983_));
 sky130_fd_sc_hd__nor2_1 _3656_ (.A(_0978_),
    .B(_0983_),
    .Y(_0371_));
 sky130_fd_sc_hd__buf_2 _3657_ (.A(_0965_),
    .X(_0984_));
 sky130_fd_sc_hd__inv_2 _3658_ (.A(\diff2[0] ),
    .Y(_0985_));
 sky130_fd_sc_hd__nor2_1 _3659_ (.A(_0984_),
    .B(_0985_),
    .Y(_0370_));
 sky130_fd_sc_hd__and2_1 _3660_ (.A(_0682_),
    .B(\diff1[36] ),
    .X(_0369_));
 sky130_fd_sc_hd__inv_2 _3661_ (.A(\diff1[35] ),
    .Y(_0986_));
 sky130_fd_sc_hd__nor2_1 _3662_ (.A(_0984_),
    .B(_0986_),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _3663_ (.A(\diff1[34] ),
    .Y(_0987_));
 sky130_fd_sc_hd__nor2_1 _3664_ (.A(_0984_),
    .B(_0987_),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_2 _3665_ (.A(\diff1[33] ),
    .Y(_0988_));
 sky130_fd_sc_hd__nor2_1 _3666_ (.A(_0984_),
    .B(_0988_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _3667_ (.A(\diff1[32] ),
    .Y(_0989_));
 sky130_fd_sc_hd__nor2_1 _3668_ (.A(_0984_),
    .B(_0989_),
    .Y(_0365_));
 sky130_fd_sc_hd__clkbuf_2 _3669_ (.A(_0965_),
    .X(_0990_));
 sky130_fd_sc_hd__inv_2 _3670_ (.A(\diff1[31] ),
    .Y(_0991_));
 sky130_fd_sc_hd__nor2_1 _3671_ (.A(_0990_),
    .B(_0991_),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_2 _3672_ (.A(\diff1[30] ),
    .Y(_0992_));
 sky130_fd_sc_hd__nor2_1 _3673_ (.A(_0990_),
    .B(_0992_),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_2 _3674_ (.A(\diff1[29] ),
    .Y(_0993_));
 sky130_fd_sc_hd__nor2_1 _3675_ (.A(_0990_),
    .B(_0993_),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _3676_ (.A(\diff1[28] ),
    .Y(_0994_));
 sky130_fd_sc_hd__nor2_1 _3677_ (.A(_0990_),
    .B(_0994_),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _3678_ (.A(\diff1[27] ),
    .Y(_0995_));
 sky130_fd_sc_hd__nor2_1 _3679_ (.A(_0990_),
    .B(_0995_),
    .Y(_0360_));
 sky130_fd_sc_hd__buf_2 _3680_ (.A(_0813_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_2 _3681_ (.A(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__inv_2 _3682_ (.A(\diff1[26] ),
    .Y(_0998_));
 sky130_fd_sc_hd__nor2_1 _3683_ (.A(_0997_),
    .B(_0998_),
    .Y(_0359_));
 sky130_fd_sc_hd__inv_2 _3684_ (.A(\diff1[25] ),
    .Y(_0999_));
 sky130_fd_sc_hd__nor2_1 _3685_ (.A(_0997_),
    .B(_0999_),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_2 _3686_ (.A(\diff1[24] ),
    .Y(_1000_));
 sky130_fd_sc_hd__nor2_1 _3687_ (.A(_0997_),
    .B(_1000_),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _3688_ (.A(\diff1[23] ),
    .Y(_1001_));
 sky130_fd_sc_hd__nor2_1 _3689_ (.A(_0997_),
    .B(_1001_),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _3690_ (.A(\diff1[22] ),
    .Y(_1002_));
 sky130_fd_sc_hd__buf_1 _3691_ (.A(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__nor2_1 _3692_ (.A(_0997_),
    .B(_1003_),
    .Y(_0355_));
 sky130_fd_sc_hd__clkbuf_2 _3693_ (.A(_0996_),
    .X(_1004_));
 sky130_fd_sc_hd__inv_2 _3694_ (.A(\diff1[21] ),
    .Y(_1005_));
 sky130_fd_sc_hd__nor2_1 _3695_ (.A(_1004_),
    .B(_1005_),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _3696_ (.A(\diff1[20] ),
    .Y(_1006_));
 sky130_fd_sc_hd__nor2_1 _3697_ (.A(_1004_),
    .B(_1006_),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _3698_ (.A(\diff1[19] ),
    .Y(_1007_));
 sky130_fd_sc_hd__nor2_1 _3699_ (.A(_1004_),
    .B(_1007_),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _3700_ (.A(\diff1[18] ),
    .Y(_1008_));
 sky130_fd_sc_hd__nor2_1 _3701_ (.A(_1004_),
    .B(_1008_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _3702_ (.A(\diff1[17] ),
    .Y(_1009_));
 sky130_fd_sc_hd__nor2_1 _3703_ (.A(_1004_),
    .B(_1009_),
    .Y(_0350_));
 sky130_fd_sc_hd__clkbuf_2 _3704_ (.A(_0996_),
    .X(_1010_));
 sky130_fd_sc_hd__inv_2 _3705_ (.A(\diff1[16] ),
    .Y(_1011_));
 sky130_fd_sc_hd__nor2_1 _3706_ (.A(_1010_),
    .B(_1011_),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _3707_ (.A(\diff1[15] ),
    .Y(_1012_));
 sky130_fd_sc_hd__nor2_1 _3708_ (.A(_1010_),
    .B(_1012_),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _3709_ (.A(\diff1[14] ),
    .Y(_1013_));
 sky130_fd_sc_hd__nor2_1 _3710_ (.A(_1010_),
    .B(_1013_),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _3711_ (.A(\diff1[13] ),
    .Y(_1014_));
 sky130_fd_sc_hd__nor2_1 _3712_ (.A(_1010_),
    .B(_1014_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _3713_ (.A(\diff1[12] ),
    .Y(_1015_));
 sky130_fd_sc_hd__nor2_1 _3714_ (.A(_1010_),
    .B(_1015_),
    .Y(_0345_));
 sky130_fd_sc_hd__clkbuf_2 _3715_ (.A(_0996_),
    .X(_1016_));
 sky130_fd_sc_hd__inv_2 _3716_ (.A(\diff1[11] ),
    .Y(_1017_));
 sky130_fd_sc_hd__nor2_1 _3717_ (.A(_1016_),
    .B(_1017_),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _3718_ (.A(\diff1[10] ),
    .Y(_1018_));
 sky130_fd_sc_hd__nor2_1 _3719_ (.A(_1016_),
    .B(_1018_),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _3720_ (.A(\diff1[9] ),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _3721_ (.A(_1016_),
    .B(_1019_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _3722_ (.A(\diff1[8] ),
    .Y(_1020_));
 sky130_fd_sc_hd__nor2_1 _3723_ (.A(_1016_),
    .B(_1020_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _3724_ (.A(\diff1[7] ),
    .Y(_1021_));
 sky130_fd_sc_hd__nor2_1 _3725_ (.A(_1016_),
    .B(_1021_),
    .Y(_0340_));
 sky130_fd_sc_hd__clkbuf_2 _3726_ (.A(_0996_),
    .X(_1022_));
 sky130_fd_sc_hd__inv_2 _3727_ (.A(\diff1[6] ),
    .Y(_1023_));
 sky130_fd_sc_hd__nor2_1 _3728_ (.A(_1022_),
    .B(_1023_),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _3729_ (.A(\diff1[5] ),
    .Y(_1024_));
 sky130_fd_sc_hd__nor2_1 _3730_ (.A(_1022_),
    .B(_1024_),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _3731_ (.A(\diff1[4] ),
    .Y(_1025_));
 sky130_fd_sc_hd__nor2_1 _3732_ (.A(_1022_),
    .B(_1025_),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _3733_ (.A(\diff1[3] ),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_1 _3734_ (.A(_1022_),
    .B(_1026_),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _3735_ (.A(\diff1[2] ),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_1 _3736_ (.A(_1022_),
    .B(_1027_),
    .Y(_0335_));
 sky130_fd_sc_hd__clkbuf_4 _3737_ (.A(_0813_),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_2 _3738_ (.A(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__inv_2 _3739_ (.A(\diff1[1] ),
    .Y(_1030_));
 sky130_fd_sc_hd__nor2_1 _3740_ (.A(_1029_),
    .B(_1030_),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _3741_ (.A(\diff1[0] ),
    .Y(_1031_));
 sky130_fd_sc_hd__nor2_1 _3742_ (.A(_1029_),
    .B(_1031_),
    .Y(_0333_));
 sky130_fd_sc_hd__a2bb2o_1 _3743_ (.A1_N(\diff2[36] ),
    .A2_N(\diff2_d[36] ),
    .B1(\diff2[36] ),
    .B2(\diff2_d[36] ),
    .X(_1032_));
 sky130_fd_sc_hd__inv_2 _3744_ (.A(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__inv_2 _3745_ (.A(\diff2_d[35] ),
    .Y(_1034_));
 sky130_fd_sc_hd__nor2_1 _3746_ (.A(\diff2[35] ),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__a21oi_2 _3747_ (.A1(\diff2[35] ),
    .A2(_1034_),
    .B1(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__inv_2 _3748_ (.A(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__a2bb2o_1 _3749_ (.A1_N(_0942_),
    .A2_N(\diff2_d[34] ),
    .B1(_0942_),
    .B2(\diff2_d[34] ),
    .X(_1038_));
 sky130_fd_sc_hd__inv_2 _3750_ (.A(\diff2_d[33] ),
    .Y(_1039_));
 sky130_fd_sc_hd__nor2_1 _3751_ (.A(\diff2[33] ),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__a21oi_2 _3752_ (.A1(\diff2[33] ),
    .A2(_1039_),
    .B1(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__inv_2 _3753_ (.A(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__a2bb2o_1 _3754_ (.A1_N(_0944_),
    .A2_N(\diff2_d[32] ),
    .B1(_0944_),
    .B2(\diff2_d[32] ),
    .X(_1043_));
 sky130_fd_sc_hd__a2bb2o_1 _3755_ (.A1_N(_0949_),
    .A2_N(\diff2_d[28] ),
    .B1(_0949_),
    .B2(\diff2_d[28] ),
    .X(_1044_));
 sky130_fd_sc_hd__inv_2 _3756_ (.A(\diff2_d[29] ),
    .Y(_1045_));
 sky130_fd_sc_hd__o22a_1 _3757_ (.A1(_0948_),
    .A2(\diff2_d[29] ),
    .B1(\diff2[29] ),
    .B2(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__inv_2 _3758_ (.A(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__or2_1 _3759_ (.A(_1044_),
    .B(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__a2bb2o_1 _3760_ (.A1_N(_0947_),
    .A2_N(\diff2_d[30] ),
    .B1(_0947_),
    .B2(\diff2_d[30] ),
    .X(_1049_));
 sky130_fd_sc_hd__inv_2 _3761_ (.A(\diff2_d[31] ),
    .Y(_1050_));
 sky130_fd_sc_hd__nor2_1 _3762_ (.A(\diff2[31] ),
    .B(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__a21oi_2 _3763_ (.A1(\diff2[31] ),
    .A2(_1050_),
    .B1(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__inv_2 _3764_ (.A(_1052_),
    .Y(_1053_));
 sky130_fd_sc_hd__or2_1 _3765_ (.A(_1049_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__or2_1 _3766_ (.A(_1048_),
    .B(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__a2bb2o_1 _3767_ (.A1_N(_0950_),
    .A2_N(\diff2_d[27] ),
    .B1(_0950_),
    .B2(\diff2_d[27] ),
    .X(_1056_));
 sky130_fd_sc_hd__a2bb2o_1 _3768_ (.A1_N(_0951_),
    .A2_N(\diff2_d[26] ),
    .B1(_0951_),
    .B2(\diff2_d[26] ),
    .X(_1057_));
 sky130_fd_sc_hd__or2_1 _3769_ (.A(_1056_),
    .B(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__inv_2 _3770_ (.A(\diff2_d[25] ),
    .Y(_1059_));
 sky130_fd_sc_hd__o22a_1 _3771_ (.A1(_0953_),
    .A2(\diff2_d[25] ),
    .B1(\diff2[25] ),
    .B2(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__inv_2 _3772_ (.A(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__a2bb2o_1 _3773_ (.A1_N(_0954_),
    .A2_N(\diff2_d[24] ),
    .B1(_0954_),
    .B2(\diff2_d[24] ),
    .X(_1062_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(_1061_),
    .B(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__or2_1 _3775_ (.A(_1058_),
    .B(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__inv_2 _3776_ (.A(\diff2_d[23] ),
    .Y(_1065_));
 sky130_fd_sc_hd__nor2_1 _3777_ (.A(\diff2[23] ),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__inv_2 _3778_ (.A(\diff2_d[21] ),
    .Y(_1067_));
 sky130_fd_sc_hd__o22a_1 _3779_ (.A1(\diff2[21] ),
    .A2(_1067_),
    .B1(_0958_),
    .B2(\diff2_d[21] ),
    .X(_1068_));
 sky130_fd_sc_hd__inv_2 _3780_ (.A(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__a2bb2o_1 _3781_ (.A1_N(_0960_),
    .A2_N(\diff2_d[20] ),
    .B1(_0960_),
    .B2(\diff2_d[20] ),
    .X(_1070_));
 sky130_fd_sc_hd__or2_1 _3782_ (.A(_1069_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__o2bb2a_1 _3783_ (.A1_N(_0961_),
    .A2_N(\diff2_d[19] ),
    .B1(_0961_),
    .B2(\diff2_d[19] ),
    .X(_1072_));
 sky130_fd_sc_hd__inv_2 _3784_ (.A(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__a2bb2o_1 _3785_ (.A1_N(_0962_),
    .A2_N(\diff2_d[18] ),
    .B1(_0962_),
    .B2(\diff2_d[18] ),
    .X(_1074_));
 sky130_fd_sc_hd__or2_1 _3786_ (.A(_1073_),
    .B(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__inv_2 _3787_ (.A(\diff2_d[17] ),
    .Y(_1076_));
 sky130_fd_sc_hd__inv_2 _3788_ (.A(\diff2_d[16] ),
    .Y(_1077_));
 sky130_fd_sc_hd__a22o_1 _3789_ (.A1(\diff2[17] ),
    .A2(_1076_),
    .B1(\diff2[16] ),
    .B2(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__o21ai_1 _3790_ (.A1(\diff2[17] ),
    .A2(_1076_),
    .B1(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__a211o_1 _3791_ (.A1(_0961_),
    .A2(\diff2_d[19] ),
    .B1(_0962_),
    .C1(\diff2_d[18] ),
    .X(_1080_));
 sky130_fd_sc_hd__o221a_1 _3792_ (.A1(_0961_),
    .A2(\diff2_d[19] ),
    .B1(_1075_),
    .B2(_1079_),
    .C1(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__or2_1 _3793_ (.A(_1071_),
    .B(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__o22ai_1 _3794_ (.A1(_0958_),
    .A2(\diff2_d[21] ),
    .B1(_0960_),
    .B2(\diff2_d[20] ),
    .Y(_1083_));
 sky130_fd_sc_hd__o21ai_1 _3795_ (.A1(\diff2[21] ),
    .A2(_1067_),
    .B1(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__a22o_1 _3796_ (.A1(_0957_),
    .A2(\diff2_d[22] ),
    .B1(_1082_),
    .B2(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__o221a_1 _3797_ (.A1(_0955_),
    .A2(\diff2_d[23] ),
    .B1(_0957_),
    .B2(\diff2_d[22] ),
    .C1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__inv_2 _3798_ (.A(\diff2_d[15] ),
    .Y(_1087_));
 sky130_fd_sc_hd__nor2_1 _3799_ (.A(\diff2[15] ),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__a21oi_2 _3800_ (.A1(\diff2[15] ),
    .A2(_1087_),
    .B1(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__inv_2 _3801_ (.A(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__a2bb2o_1 _3802_ (.A1_N(_0968_),
    .A2_N(\diff2_d[14] ),
    .B1(_0968_),
    .B2(\diff2_d[14] ),
    .X(_1091_));
 sky130_fd_sc_hd__or2_1 _3803_ (.A(_1090_),
    .B(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__inv_2 _3804_ (.A(\diff2_d[13] ),
    .Y(_1093_));
 sky130_fd_sc_hd__o22a_1 _3805_ (.A1(_0969_),
    .A2(\diff2_d[13] ),
    .B1(\diff2[13] ),
    .B2(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__inv_2 _3806_ (.A(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__a2bb2o_1 _3807_ (.A1_N(_0970_),
    .A2_N(\diff2_d[12] ),
    .B1(_0970_),
    .B2(\diff2_d[12] ),
    .X(_1096_));
 sky130_fd_sc_hd__or2_1 _3808_ (.A(_1095_),
    .B(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__or2_1 _3809_ (.A(_1092_),
    .B(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__a2bb2o_1 _3810_ (.A1_N(_0971_),
    .A2_N(\diff2_d[11] ),
    .B1(_0971_),
    .B2(\diff2_d[11] ),
    .X(_1099_));
 sky130_fd_sc_hd__a2bb2o_1 _3811_ (.A1_N(_0973_),
    .A2_N(\diff2_d[10] ),
    .B1(_0973_),
    .B2(\diff2_d[10] ),
    .X(_1100_));
 sky130_fd_sc_hd__or2_1 _3812_ (.A(_1099_),
    .B(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__inv_2 _3813_ (.A(\diff2_d[9] ),
    .Y(_1102_));
 sky130_fd_sc_hd__o22a_1 _3814_ (.A1(_0974_),
    .A2(\diff2_d[9] ),
    .B1(\diff2[9] ),
    .B2(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__inv_2 _3815_ (.A(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__a2bb2o_1 _3816_ (.A1_N(_0975_),
    .A2_N(\diff2_d[8] ),
    .B1(_0975_),
    .B2(\diff2_d[8] ),
    .X(_1105_));
 sky130_fd_sc_hd__or2_1 _3817_ (.A(_1104_),
    .B(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__or2_1 _3818_ (.A(_1101_),
    .B(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__inv_2 _3819_ (.A(\diff2_d[7] ),
    .Y(_1108_));
 sky130_fd_sc_hd__nor2_1 _3820_ (.A(\diff2[7] ),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__a21oi_2 _3821_ (.A1(\diff2[7] ),
    .A2(_1108_),
    .B1(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__inv_2 _3822_ (.A(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__a2bb2o_1 _3823_ (.A1_N(_0977_),
    .A2_N(\diff2_d[6] ),
    .B1(_0977_),
    .B2(\diff2_d[6] ),
    .X(_1112_));
 sky130_fd_sc_hd__nor2_1 _3824_ (.A(_0979_),
    .B(\diff2_d[5] ),
    .Y(_1113_));
 sky130_fd_sc_hd__nor2_4 _3825_ (.A(_0980_),
    .B(\diff2_d[4] ),
    .Y(_1114_));
 sky130_fd_sc_hd__o2bb2a_1 _3826_ (.A1_N(_0979_),
    .A2_N(\diff2_d[5] ),
    .B1(_1113_),
    .B2(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__inv_2 _3827_ (.A(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__o32a_1 _3828_ (.A1(_0977_),
    .A2(\diff2_d[6] ),
    .A3(_1109_),
    .B1(_0976_),
    .B2(\diff2_d[7] ),
    .X(_1117_));
 sky130_fd_sc_hd__a21oi_2 _3829_ (.A1(_0979_),
    .A2(\diff2_d[5] ),
    .B1(_1113_),
    .Y(_1118_));
 sky130_fd_sc_hd__a21oi_4 _3830_ (.A1(_0980_),
    .A2(\diff2_d[4] ),
    .B1(_1114_),
    .Y(_1119_));
 sky130_fd_sc_hd__nand2_1 _3831_ (.A(_1118_),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__inv_2 _3832_ (.A(\diff2_d[3] ),
    .Y(_1121_));
 sky130_fd_sc_hd__nor2_1 _3833_ (.A(\diff2[3] ),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__a21oi_2 _3834_ (.A1(\diff2[3] ),
    .A2(_1121_),
    .B1(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__inv_2 _3835_ (.A(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__a2bb2o_1 _3836_ (.A1_N(_0982_),
    .A2_N(\diff2_d[2] ),
    .B1(_0982_),
    .B2(\diff2_d[2] ),
    .X(_1125_));
 sky130_fd_sc_hd__inv_2 _3837_ (.A(\diff2_d[0] ),
    .Y(_1126_));
 sky130_fd_sc_hd__inv_2 _3838_ (.A(\diff2_d[1] ),
    .Y(_1127_));
 sky130_fd_sc_hd__o22a_1 _3839_ (.A1(_0983_),
    .A2(\diff2_d[1] ),
    .B1(\diff2[1] ),
    .B2(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__o21ai_1 _3840_ (.A1(\diff2[0] ),
    .A2(_1126_),
    .B1(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__o21ai_2 _3841_ (.A1(_0983_),
    .A2(\diff2_d[1] ),
    .B1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__inv_2 _3842_ (.A(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__o32a_1 _3843_ (.A1(_0982_),
    .A2(\diff2_d[2] ),
    .A3(_1122_),
    .B1(_0981_),
    .B2(\diff2_d[3] ),
    .X(_1132_));
 sky130_fd_sc_hd__o31a_1 _3844_ (.A1(_1124_),
    .A2(_1125_),
    .A3(_1131_),
    .B1(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__or4_4 _3845_ (.A(_1111_),
    .B(_1112_),
    .C(_1120_),
    .D(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__o311a_2 _3846_ (.A1(_1111_),
    .A2(_1112_),
    .A3(_1116_),
    .B1(_1117_),
    .C1(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__o22ai_1 _3847_ (.A1(_0969_),
    .A2(\diff2_d[13] ),
    .B1(_0970_),
    .B2(\diff2_d[12] ),
    .Y(_1136_));
 sky130_fd_sc_hd__o21ai_1 _3848_ (.A1(\diff2[13] ),
    .A2(_1093_),
    .B1(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__o22ai_1 _3849_ (.A1(_0974_),
    .A2(\diff2_d[9] ),
    .B1(_0975_),
    .B2(\diff2_d[8] ),
    .Y(_1138_));
 sky130_fd_sc_hd__o21ai_1 _3850_ (.A1(\diff2[9] ),
    .A2(_1102_),
    .B1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__a211o_1 _3851_ (.A1(_0971_),
    .A2(\diff2_d[11] ),
    .B1(_0973_),
    .C1(\diff2_d[10] ),
    .X(_1140_));
 sky130_fd_sc_hd__o221a_1 _3852_ (.A1(_0971_),
    .A2(\diff2_d[11] ),
    .B1(_1101_),
    .B2(_1139_),
    .C1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__o32a_1 _3853_ (.A1(_0968_),
    .A2(\diff2_d[14] ),
    .A3(_1088_),
    .B1(_0967_),
    .B2(\diff2_d[15] ),
    .X(_1142_));
 sky130_fd_sc_hd__o221a_1 _3854_ (.A1(_1092_),
    .A2(_1137_),
    .B1(_1098_),
    .B2(_1141_),
    .C1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__o31a_2 _3855_ (.A1(_1098_),
    .A2(_1107_),
    .A3(_1135_),
    .B1(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__o22a_1 _3856_ (.A1(\diff2[17] ),
    .A2(_1076_),
    .B1(_0963_),
    .B2(\diff2_d[17] ),
    .X(_1145_));
 sky130_fd_sc_hd__inv_2 _3857_ (.A(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__o22a_1 _3858_ (.A1(_0964_),
    .A2(\diff2_d[16] ),
    .B1(\diff2[16] ),
    .B2(_1077_),
    .X(_1147_));
 sky130_fd_sc_hd__inv_2 _3859_ (.A(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__or2_1 _3860_ (.A(_1146_),
    .B(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__or2_1 _3861_ (.A(_1075_),
    .B(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__a21oi_2 _3862_ (.A1(\diff2[23] ),
    .A2(_1065_),
    .B1(_1066_),
    .Y(_1151_));
 sky130_fd_sc_hd__inv_2 _3863_ (.A(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__o2bb2a_1 _3864_ (.A1_N(_0957_),
    .A2_N(\diff2_d[22] ),
    .B1(_0956_),
    .B2(\diff2_d[22] ),
    .X(_1153_));
 sky130_fd_sc_hd__or4b_4 _3865_ (.A(_1150_),
    .B(_1152_),
    .C(_1071_),
    .D_N(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__o22a_2 _3866_ (.A1(_1066_),
    .A2(_1086_),
    .B1(_1144_),
    .B2(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__a2bb2o_1 _3867_ (.A1_N(_0949_),
    .A2_N(\diff2_d[28] ),
    .B1(\diff2[29] ),
    .B2(_1045_),
    .X(_1156_));
 sky130_fd_sc_hd__o21ai_1 _3868_ (.A1(\diff2[29] ),
    .A2(_1045_),
    .B1(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__o22ai_1 _3869_ (.A1(_0953_),
    .A2(\diff2_d[25] ),
    .B1(_0954_),
    .B2(\diff2_d[24] ),
    .Y(_1158_));
 sky130_fd_sc_hd__o21ai_1 _3870_ (.A1(\diff2[25] ),
    .A2(_1059_),
    .B1(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__a211o_1 _3871_ (.A1(_0950_),
    .A2(\diff2_d[27] ),
    .B1(_0951_),
    .C1(\diff2_d[26] ),
    .X(_1160_));
 sky130_fd_sc_hd__o221a_1 _3872_ (.A1(_0950_),
    .A2(\diff2_d[27] ),
    .B1(_1058_),
    .B2(_1159_),
    .C1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__o32a_1 _3873_ (.A1(_0947_),
    .A2(\diff2_d[30] ),
    .A3(_1051_),
    .B1(_0945_),
    .B2(\diff2_d[31] ),
    .X(_1162_));
 sky130_fd_sc_hd__o221a_1 _3874_ (.A1(_1054_),
    .A2(_1157_),
    .B1(_1055_),
    .B2(_1161_),
    .C1(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__o31a_1 _3875_ (.A1(_1055_),
    .A2(_1064_),
    .A3(_1155_),
    .B1(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__o32a_1 _3876_ (.A1(_0944_),
    .A2(\diff2_d[32] ),
    .A3(_1040_),
    .B1(_0943_),
    .B2(\diff2_d[33] ),
    .X(_1165_));
 sky130_fd_sc_hd__o31a_1 _3877_ (.A1(_1042_),
    .A2(_1043_),
    .A3(_1164_),
    .B1(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__o32a_1 _3878_ (.A1(_0942_),
    .A2(\diff2_d[34] ),
    .A3(_1035_),
    .B1(_0941_),
    .B2(\diff2_d[35] ),
    .X(_1167_));
 sky130_fd_sc_hd__o31a_1 _3879_ (.A1(_1037_),
    .A2(_1038_),
    .A3(_1166_),
    .B1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__inv_2 _3880_ (.A(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__o221a_1 _3881_ (.A1(_1033_),
    .A2(_1168_),
    .B1(_1032_),
    .B2(_1169_),
    .C1(_0812_),
    .X(_0332_));
 sky130_fd_sc_hd__or2_1 _3882_ (.A(_1166_),
    .B(_1038_),
    .X(_1170_));
 sky130_fd_sc_hd__o21ai_1 _3883_ (.A1(_0942_),
    .A2(\diff2_d[34] ),
    .B1(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__inv_2 _3884_ (.A(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__o221a_1 _3885_ (.A1(_1037_),
    .A2(_1172_),
    .B1(_1036_),
    .B2(_1171_),
    .C1(_0812_),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_2 _3886_ (.A(_0681_),
    .X(_1173_));
 sky130_fd_sc_hd__nand2_1 _3887_ (.A(_1166_),
    .B(_1038_),
    .Y(_1174_));
 sky130_fd_sc_hd__and3_1 _3888_ (.A(_1173_),
    .B(_1170_),
    .C(_1174_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_1 _3889_ (.A(_1164_),
    .B(_1043_),
    .X(_1175_));
 sky130_fd_sc_hd__o21ai_1 _3890_ (.A1(_0944_),
    .A2(\diff2_d[32] ),
    .B1(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__inv_2 _3891_ (.A(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__o221a_1 _3892_ (.A1(_1042_),
    .A2(_1177_),
    .B1(_1041_),
    .B2(_1176_),
    .C1(_0812_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _3893_ (.A(_1164_),
    .B(_1043_),
    .Y(_1178_));
 sky130_fd_sc_hd__and3_1 _3894_ (.A(_1173_),
    .B(_1175_),
    .C(_1178_),
    .X(_0328_));
 sky130_fd_sc_hd__inv_2 _3895_ (.A(_1049_),
    .Y(_1179_));
 sky130_fd_sc_hd__o21ai_2 _3896_ (.A1(_1155_),
    .A2(_1064_),
    .B1(_1161_),
    .Y(_1180_));
 sky130_fd_sc_hd__inv_2 _3897_ (.A(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__o21ai_1 _3898_ (.A1(_1048_),
    .A2(_1181_),
    .B1(_1157_),
    .Y(_1182_));
 sky130_fd_sc_hd__nand2_1 _3899_ (.A(_1179_),
    .B(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__o21ai_1 _3900_ (.A1(_0947_),
    .A2(\diff2_d[30] ),
    .B1(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__inv_2 _3901_ (.A(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__clkbuf_2 _3902_ (.A(_0705_),
    .X(_1186_));
 sky130_fd_sc_hd__o221a_1 _3903_ (.A1(_1053_),
    .A2(_1185_),
    .B1(_1052_),
    .B2(_1184_),
    .C1(_1186_),
    .X(_0327_));
 sky130_fd_sc_hd__o211a_1 _3904_ (.A1(_1179_),
    .A2(_1182_),
    .B1(_0849_),
    .C1(_1183_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _3905_ (.A(_1044_),
    .B(_1181_),
    .X(_1187_));
 sky130_fd_sc_hd__o21ai_1 _3906_ (.A1(_0949_),
    .A2(\diff2_d[28] ),
    .B1(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__inv_2 _3907_ (.A(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__o221a_1 _3908_ (.A1(_1047_),
    .A2(_1189_),
    .B1(_1046_),
    .B2(_1188_),
    .C1(_1186_),
    .X(_0325_));
 sky130_fd_sc_hd__inv_2 _3909_ (.A(_1044_),
    .Y(_1190_));
 sky130_fd_sc_hd__o211a_1 _3910_ (.A1(_1190_),
    .A2(_1180_),
    .B1(_0849_),
    .C1(_1187_),
    .X(_0324_));
 sky130_fd_sc_hd__inv_2 _3911_ (.A(_1057_),
    .Y(_1191_));
 sky130_fd_sc_hd__o21ai_1 _3912_ (.A1(_1155_),
    .A2(_1063_),
    .B1(_1159_),
    .Y(_1192_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(_1191_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__o21ai_1 _3914_ (.A1(_0951_),
    .A2(\diff2_d[26] ),
    .B1(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__inv_2 _3915_ (.A(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__inv_2 _3916_ (.A(_1056_),
    .Y(_1196_));
 sky130_fd_sc_hd__o221a_1 _3917_ (.A1(_1056_),
    .A2(_1195_),
    .B1(_1196_),
    .B2(_1194_),
    .C1(_1186_),
    .X(_0323_));
 sky130_fd_sc_hd__o211a_1 _3918_ (.A1(_1191_),
    .A2(_1192_),
    .B1(_0849_),
    .C1(_1193_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _3919_ (.A(_1155_),
    .B(_1062_),
    .X(_1197_));
 sky130_fd_sc_hd__o21ai_1 _3920_ (.A1(_0954_),
    .A2(\diff2_d[24] ),
    .B1(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__inv_2 _3921_ (.A(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__o221a_1 _3922_ (.A1(_1061_),
    .A2(_1199_),
    .B1(_1060_),
    .B2(_1198_),
    .C1(_1186_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2_1 _3923_ (.A(_1155_),
    .B(_1062_),
    .Y(_1200_));
 sky130_fd_sc_hd__and3_1 _3924_ (.A(_1173_),
    .B(_1197_),
    .C(_1200_),
    .X(_0320_));
 sky130_fd_sc_hd__o21ai_1 _3925_ (.A1(_1144_),
    .A2(_1150_),
    .B1(_1081_),
    .Y(_1201_));
 sky130_fd_sc_hd__inv_2 _3926_ (.A(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__o21ai_1 _3927_ (.A1(_1071_),
    .A2(_1202_),
    .B1(_1084_),
    .Y(_1203_));
 sky130_fd_sc_hd__nand2_1 _3928_ (.A(_1153_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__o21ai_1 _3929_ (.A1(_0957_),
    .A2(\diff2_d[22] ),
    .B1(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__inv_2 _3930_ (.A(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__o221a_1 _3931_ (.A1(_1152_),
    .A2(_1206_),
    .B1(_1151_),
    .B2(_1205_),
    .C1(_1186_),
    .X(_0319_));
 sky130_fd_sc_hd__o211a_1 _3932_ (.A1(_1153_),
    .A2(_1203_),
    .B1(_0849_),
    .C1(_1204_),
    .X(_0318_));
 sky130_fd_sc_hd__or2_1 _3933_ (.A(_1070_),
    .B(_1202_),
    .X(_1207_));
 sky130_fd_sc_hd__o21ai_1 _3934_ (.A1(_0960_),
    .A2(\diff2_d[20] ),
    .B1(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__inv_2 _3935_ (.A(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__clkbuf_2 _3936_ (.A(_0705_),
    .X(_1210_));
 sky130_fd_sc_hd__o221a_1 _3937_ (.A1(_1069_),
    .A2(_1209_),
    .B1(_1068_),
    .B2(_1208_),
    .C1(_1210_),
    .X(_0317_));
 sky130_fd_sc_hd__inv_2 _3938_ (.A(_1070_),
    .Y(_1211_));
 sky130_fd_sc_hd__clkbuf_2 _3939_ (.A(_0830_),
    .X(_1212_));
 sky130_fd_sc_hd__o211a_1 _3940_ (.A1(_1211_),
    .A2(_1201_),
    .B1(_1212_),
    .C1(_1207_),
    .X(_0316_));
 sky130_fd_sc_hd__inv_2 _3941_ (.A(_1074_),
    .Y(_1213_));
 sky130_fd_sc_hd__o21ai_1 _3942_ (.A1(_1144_),
    .A2(_1149_),
    .B1(_1079_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _3943_ (.A(_1213_),
    .B(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__o21ai_1 _3944_ (.A1(_0962_),
    .A2(\diff2_d[18] ),
    .B1(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__inv_2 _3945_ (.A(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__o221a_1 _3946_ (.A1(_1073_),
    .A2(_1217_),
    .B1(_1072_),
    .B2(_1216_),
    .C1(_1210_),
    .X(_0315_));
 sky130_fd_sc_hd__o211a_1 _3947_ (.A1(_1213_),
    .A2(_1214_),
    .B1(_1212_),
    .C1(_1215_),
    .X(_0314_));
 sky130_fd_sc_hd__or2_1 _3948_ (.A(_1144_),
    .B(_1148_),
    .X(_1218_));
 sky130_fd_sc_hd__o21ai_1 _3949_ (.A1(_0964_),
    .A2(\diff2_d[16] ),
    .B1(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__inv_2 _3950_ (.A(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__o221a_1 _3951_ (.A1(_1146_),
    .A2(_1220_),
    .B1(_1145_),
    .B2(_1219_),
    .C1(_1210_),
    .X(_0313_));
 sky130_fd_sc_hd__inv_2 _3952_ (.A(_1144_),
    .Y(_1221_));
 sky130_fd_sc_hd__o211a_1 _3953_ (.A1(_1221_),
    .A2(_1147_),
    .B1(_1212_),
    .C1(_1218_),
    .X(_0312_));
 sky130_fd_sc_hd__inv_2 _3954_ (.A(_1091_),
    .Y(_1222_));
 sky130_fd_sc_hd__o21ai_1 _3955_ (.A1(_1135_),
    .A2(_1107_),
    .B1(_1141_),
    .Y(_1223_));
 sky130_fd_sc_hd__inv_2 _3956_ (.A(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__o21ai_1 _3957_ (.A1(_1097_),
    .A2(_1224_),
    .B1(_1137_),
    .Y(_1225_));
 sky130_fd_sc_hd__nand2_1 _3958_ (.A(_1222_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__o21ai_1 _3959_ (.A1(_0968_),
    .A2(\diff2_d[14] ),
    .B1(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__inv_2 _3960_ (.A(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__o221a_1 _3961_ (.A1(_1090_),
    .A2(_1228_),
    .B1(_1089_),
    .B2(_1227_),
    .C1(_1210_),
    .X(_0311_));
 sky130_fd_sc_hd__o211a_1 _3962_ (.A1(_1222_),
    .A2(_1225_),
    .B1(_1212_),
    .C1(_1226_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _3963_ (.A(_1096_),
    .B(_1224_),
    .X(_1229_));
 sky130_fd_sc_hd__o21ai_1 _3964_ (.A1(_0970_),
    .A2(\diff2_d[12] ),
    .B1(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__inv_2 _3965_ (.A(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__o221a_1 _3966_ (.A1(_1095_),
    .A2(_1231_),
    .B1(_1094_),
    .B2(_1230_),
    .C1(_1210_),
    .X(_0309_));
 sky130_fd_sc_hd__inv_2 _3967_ (.A(_1096_),
    .Y(_1232_));
 sky130_fd_sc_hd__o211a_1 _3968_ (.A1(_1232_),
    .A2(_1223_),
    .B1(_1212_),
    .C1(_1229_),
    .X(_0308_));
 sky130_fd_sc_hd__inv_2 _3969_ (.A(_1100_),
    .Y(_1233_));
 sky130_fd_sc_hd__o21ai_1 _3970_ (.A1(_1135_),
    .A2(_1106_),
    .B1(_1139_),
    .Y(_1234_));
 sky130_fd_sc_hd__nand2_1 _3971_ (.A(_1233_),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__o21ai_1 _3972_ (.A1(_0973_),
    .A2(\diff2_d[10] ),
    .B1(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__inv_2 _3973_ (.A(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__inv_2 _3974_ (.A(_1099_),
    .Y(_1238_));
 sky130_fd_sc_hd__clkbuf_2 _3975_ (.A(_0680_),
    .X(_1239_));
 sky130_fd_sc_hd__buf_2 _3976_ (.A(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__o221a_1 _3977_ (.A1(_1099_),
    .A2(_1237_),
    .B1(_1238_),
    .B2(_1236_),
    .C1(_1240_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_2 _3978_ (.A(_0830_),
    .X(_1241_));
 sky130_fd_sc_hd__o211a_1 _3979_ (.A1(_1233_),
    .A2(_1234_),
    .B1(_1241_),
    .C1(_1235_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _3980_ (.A(_1135_),
    .B(_1105_),
    .X(_1242_));
 sky130_fd_sc_hd__o21ai_1 _3981_ (.A1(_0975_),
    .A2(\diff2_d[8] ),
    .B1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__inv_2 _3982_ (.A(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__o221a_1 _3983_ (.A1(_1104_),
    .A2(_1244_),
    .B1(_1103_),
    .B2(_1243_),
    .C1(_1240_),
    .X(_0305_));
 sky130_fd_sc_hd__nand2_1 _3984_ (.A(_1135_),
    .B(_1105_),
    .Y(_1245_));
 sky130_fd_sc_hd__and3_1 _3985_ (.A(_1173_),
    .B(_1242_),
    .C(_1245_),
    .X(_0304_));
 sky130_fd_sc_hd__inv_2 _3986_ (.A(_1112_),
    .Y(_1246_));
 sky130_fd_sc_hd__inv_2 _3987_ (.A(_1133_),
    .Y(_1247_));
 sky130_fd_sc_hd__a31o_1 _3988_ (.A1(_1118_),
    .A2(_1119_),
    .A3(_1247_),
    .B1(_1115_),
    .X(_1248_));
 sky130_fd_sc_hd__nand2_1 _3989_ (.A(_1246_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__o21ai_1 _3990_ (.A1(_0977_),
    .A2(\diff2_d[6] ),
    .B1(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__inv_2 _3991_ (.A(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__o221a_1 _3992_ (.A1(_1111_),
    .A2(_1251_),
    .B1(_1110_),
    .B2(_1250_),
    .C1(_1240_),
    .X(_0303_));
 sky130_fd_sc_hd__o211a_1 _3993_ (.A1(_1246_),
    .A2(_1248_),
    .B1(_1241_),
    .C1(_1249_),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _3994_ (.A(_1247_),
    .B(_1119_),
    .Y(_1252_));
 sky130_fd_sc_hd__inv_2 _3995_ (.A(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__buf_2 _3996_ (.A(_0681_),
    .X(_1254_));
 sky130_fd_sc_hd__o21ai_1 _3997_ (.A1(_1114_),
    .A2(_1253_),
    .B1(_1118_),
    .Y(_1255_));
 sky130_fd_sc_hd__o311a_1 _3998_ (.A1(_1114_),
    .A2(_1253_),
    .A3(_1118_),
    .B1(_1254_),
    .C1(_1255_),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_1 _3999_ (.A1(_1247_),
    .A2(_1119_),
    .B1(_1241_),
    .C1(_1252_),
    .X(_0300_));
 sky130_fd_sc_hd__or2_1 _4000_ (.A(_1131_),
    .B(_1125_),
    .X(_1256_));
 sky130_fd_sc_hd__o21ai_1 _4001_ (.A1(_0982_),
    .A2(\diff2_d[2] ),
    .B1(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__inv_2 _4002_ (.A(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__o221a_1 _4003_ (.A1(_1124_),
    .A2(_1258_),
    .B1(_1123_),
    .B2(_1257_),
    .C1(_1240_),
    .X(_0299_));
 sky130_fd_sc_hd__inv_2 _4004_ (.A(_1125_),
    .Y(_1259_));
 sky130_fd_sc_hd__o211a_1 _4005_ (.A1(_1130_),
    .A2(_1259_),
    .B1(_1241_),
    .C1(_1256_),
    .X(_0298_));
 sky130_fd_sc_hd__o311a_1 _4006_ (.A1(\diff2[0] ),
    .A2(_1126_),
    .A3(_1128_),
    .B1(_1254_),
    .C1(_1129_),
    .X(_0297_));
 sky130_fd_sc_hd__o22a_1 _4007_ (.A1(\diff2[0] ),
    .A2(_1126_),
    .B1(_0985_),
    .B2(\diff2_d[0] ),
    .X(_1260_));
 sky130_fd_sc_hd__nor2_1 _4008_ (.A(_1029_),
    .B(_1260_),
    .Y(_0296_));
 sky130_fd_sc_hd__a2bb2o_1 _4009_ (.A1_N(\diff1[36] ),
    .A2_N(\diff1_d[36] ),
    .B1(\diff1[36] ),
    .B2(\diff1_d[36] ),
    .X(_1261_));
 sky130_fd_sc_hd__inv_2 _4010_ (.A(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__inv_2 _4011_ (.A(\diff1_d[35] ),
    .Y(_1263_));
 sky130_fd_sc_hd__nor2_1 _4012_ (.A(\diff1[35] ),
    .B(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__a21oi_2 _4013_ (.A1(\diff1[35] ),
    .A2(_1263_),
    .B1(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__inv_2 _4014_ (.A(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__a2bb2o_1 _4015_ (.A1_N(_0987_),
    .A2_N(\diff1_d[34] ),
    .B1(_0987_),
    .B2(\diff1_d[34] ),
    .X(_1267_));
 sky130_fd_sc_hd__inv_2 _4016_ (.A(\diff1_d[33] ),
    .Y(_1268_));
 sky130_fd_sc_hd__nor2_1 _4017_ (.A(\diff1[33] ),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__a21oi_2 _4018_ (.A1(\diff1[33] ),
    .A2(_1268_),
    .B1(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__inv_2 _4019_ (.A(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__a2bb2o_1 _4020_ (.A1_N(_0989_),
    .A2_N(\diff1_d[32] ),
    .B1(_0989_),
    .B2(\diff1_d[32] ),
    .X(_1272_));
 sky130_fd_sc_hd__a2bb2o_1 _4021_ (.A1_N(_0994_),
    .A2_N(\diff1_d[28] ),
    .B1(_0994_),
    .B2(\diff1_d[28] ),
    .X(_1273_));
 sky130_fd_sc_hd__inv_2 _4022_ (.A(\diff1_d[29] ),
    .Y(_1274_));
 sky130_fd_sc_hd__o22a_1 _4023_ (.A1(_0993_),
    .A2(\diff1_d[29] ),
    .B1(\diff1[29] ),
    .B2(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__inv_2 _4024_ (.A(_1275_),
    .Y(_1276_));
 sky130_fd_sc_hd__or2_1 _4025_ (.A(_1273_),
    .B(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__a2bb2o_1 _4026_ (.A1_N(_0992_),
    .A2_N(\diff1_d[30] ),
    .B1(_0992_),
    .B2(\diff1_d[30] ),
    .X(_1278_));
 sky130_fd_sc_hd__inv_2 _4027_ (.A(\diff1_d[31] ),
    .Y(_1279_));
 sky130_fd_sc_hd__nor2_1 _4028_ (.A(\diff1[31] ),
    .B(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__a21oi_2 _4029_ (.A1(\diff1[31] ),
    .A2(_1279_),
    .B1(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__inv_2 _4030_ (.A(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__or2_1 _4031_ (.A(_1278_),
    .B(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__or2_1 _4032_ (.A(_1277_),
    .B(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a2bb2o_1 _4033_ (.A1_N(_0995_),
    .A2_N(\diff1_d[27] ),
    .B1(_0995_),
    .B2(\diff1_d[27] ),
    .X(_1285_));
 sky130_fd_sc_hd__a2bb2o_1 _4034_ (.A1_N(_0998_),
    .A2_N(\diff1_d[26] ),
    .B1(_0998_),
    .B2(\diff1_d[26] ),
    .X(_1286_));
 sky130_fd_sc_hd__or2_1 _4035_ (.A(_1285_),
    .B(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__inv_2 _4036_ (.A(\diff1_d[25] ),
    .Y(_1288_));
 sky130_fd_sc_hd__o22a_1 _4037_ (.A1(_0999_),
    .A2(\diff1_d[25] ),
    .B1(\diff1[25] ),
    .B2(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__inv_2 _4038_ (.A(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__a2bb2o_1 _4039_ (.A1_N(_1000_),
    .A2_N(\diff1_d[24] ),
    .B1(_1000_),
    .B2(\diff1_d[24] ),
    .X(_1291_));
 sky130_fd_sc_hd__or2_1 _4040_ (.A(_1290_),
    .B(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__or2_1 _4041_ (.A(_1287_),
    .B(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__inv_2 _4042_ (.A(\diff1_d[23] ),
    .Y(_1294_));
 sky130_fd_sc_hd__nor2_1 _4043_ (.A(\diff1[23] ),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_2 _4044_ (.A(\diff1_d[21] ),
    .Y(_1296_));
 sky130_fd_sc_hd__o22a_1 _4045_ (.A1(\diff1[21] ),
    .A2(_1296_),
    .B1(_1005_),
    .B2(\diff1_d[21] ),
    .X(_1297_));
 sky130_fd_sc_hd__inv_2 _4046_ (.A(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__a2bb2o_1 _4047_ (.A1_N(_1006_),
    .A2_N(\diff1_d[20] ),
    .B1(_1006_),
    .B2(\diff1_d[20] ),
    .X(_1299_));
 sky130_fd_sc_hd__or2_1 _4048_ (.A(_1298_),
    .B(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__o2bb2a_1 _4049_ (.A1_N(_1007_),
    .A2_N(\diff1_d[19] ),
    .B1(_1007_),
    .B2(\diff1_d[19] ),
    .X(_1301_));
 sky130_fd_sc_hd__inv_2 _4050_ (.A(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__a2bb2o_1 _4051_ (.A1_N(_1008_),
    .A2_N(\diff1_d[18] ),
    .B1(_1008_),
    .B2(\diff1_d[18] ),
    .X(_1303_));
 sky130_fd_sc_hd__or2_1 _4052_ (.A(_1302_),
    .B(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__inv_2 _4053_ (.A(\diff1_d[17] ),
    .Y(_1305_));
 sky130_fd_sc_hd__inv_2 _4054_ (.A(\diff1_d[16] ),
    .Y(_1306_));
 sky130_fd_sc_hd__a22o_1 _4055_ (.A1(\diff1[17] ),
    .A2(_1305_),
    .B1(\diff1[16] ),
    .B2(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__o21ai_1 _4056_ (.A1(\diff1[17] ),
    .A2(_1305_),
    .B1(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__a211o_1 _4057_ (.A1(_1007_),
    .A2(\diff1_d[19] ),
    .B1(_1008_),
    .C1(\diff1_d[18] ),
    .X(_1309_));
 sky130_fd_sc_hd__o221a_1 _4058_ (.A1(_1007_),
    .A2(\diff1_d[19] ),
    .B1(_1304_),
    .B2(_1308_),
    .C1(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__or2_1 _4059_ (.A(_1300_),
    .B(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__o22ai_1 _4060_ (.A1(_1005_),
    .A2(\diff1_d[21] ),
    .B1(_1006_),
    .B2(\diff1_d[20] ),
    .Y(_1312_));
 sky130_fd_sc_hd__o21ai_1 _4061_ (.A1(\diff1[21] ),
    .A2(_1296_),
    .B1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__a22o_1 _4062_ (.A1(_1003_),
    .A2(\diff1_d[22] ),
    .B1(_1311_),
    .B2(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__o221a_1 _4063_ (.A1(_1001_),
    .A2(\diff1_d[23] ),
    .B1(_1003_),
    .B2(\diff1_d[22] ),
    .C1(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__inv_2 _4064_ (.A(\diff1_d[15] ),
    .Y(_1316_));
 sky130_fd_sc_hd__nor2_1 _4065_ (.A(\diff1[15] ),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__a21oi_2 _4066_ (.A1(\diff1[15] ),
    .A2(_1316_),
    .B1(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__inv_2 _4067_ (.A(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__a2bb2o_1 _4068_ (.A1_N(_1013_),
    .A2_N(\diff1_d[14] ),
    .B1(_1013_),
    .B2(\diff1_d[14] ),
    .X(_1320_));
 sky130_fd_sc_hd__or2_1 _4069_ (.A(_1319_),
    .B(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__inv_2 _4070_ (.A(\diff1_d[13] ),
    .Y(_1322_));
 sky130_fd_sc_hd__o22a_1 _4071_ (.A1(_1014_),
    .A2(\diff1_d[13] ),
    .B1(\diff1[13] ),
    .B2(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__inv_2 _4072_ (.A(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__a2bb2o_1 _4073_ (.A1_N(_1015_),
    .A2_N(\diff1_d[12] ),
    .B1(_1015_),
    .B2(\diff1_d[12] ),
    .X(_1325_));
 sky130_fd_sc_hd__or2_1 _4074_ (.A(_1324_),
    .B(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__or2_1 _4075_ (.A(_1321_),
    .B(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__a2bb2o_1 _4076_ (.A1_N(_1017_),
    .A2_N(\diff1_d[11] ),
    .B1(_1017_),
    .B2(\diff1_d[11] ),
    .X(_1328_));
 sky130_fd_sc_hd__a2bb2o_1 _4077_ (.A1_N(_1018_),
    .A2_N(\diff1_d[10] ),
    .B1(_1018_),
    .B2(\diff1_d[10] ),
    .X(_1329_));
 sky130_fd_sc_hd__or2_1 _4078_ (.A(_1328_),
    .B(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__inv_2 _4079_ (.A(\diff1_d[9] ),
    .Y(_1331_));
 sky130_fd_sc_hd__o22a_1 _4080_ (.A1(_1019_),
    .A2(\diff1_d[9] ),
    .B1(\diff1[9] ),
    .B2(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__inv_2 _4081_ (.A(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__a2bb2o_1 _4082_ (.A1_N(_1020_),
    .A2_N(\diff1_d[8] ),
    .B1(_1020_),
    .B2(\diff1_d[8] ),
    .X(_1334_));
 sky130_fd_sc_hd__or2_1 _4083_ (.A(_1333_),
    .B(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__or2_1 _4084_ (.A(_1330_),
    .B(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__inv_2 _4085_ (.A(\diff1_d[7] ),
    .Y(_1337_));
 sky130_fd_sc_hd__nor2_1 _4086_ (.A(\diff1[7] ),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__a21oi_2 _4087_ (.A1(\diff1[7] ),
    .A2(_1337_),
    .B1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__inv_2 _4088_ (.A(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__a2bb2o_1 _4089_ (.A1_N(_1023_),
    .A2_N(\diff1_d[6] ),
    .B1(_1023_),
    .B2(\diff1_d[6] ),
    .X(_1341_));
 sky130_fd_sc_hd__nor2_1 _4090_ (.A(_1024_),
    .B(\diff1_d[5] ),
    .Y(_1342_));
 sky130_fd_sc_hd__nor2_4 _4091_ (.A(_1025_),
    .B(\diff1_d[4] ),
    .Y(_1343_));
 sky130_fd_sc_hd__o2bb2a_1 _4092_ (.A1_N(_1024_),
    .A2_N(\diff1_d[5] ),
    .B1(_1342_),
    .B2(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__inv_2 _4093_ (.A(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__o32a_1 _4094_ (.A1(_1023_),
    .A2(\diff1_d[6] ),
    .A3(_1338_),
    .B1(_1021_),
    .B2(\diff1_d[7] ),
    .X(_1346_));
 sky130_fd_sc_hd__a21oi_2 _4095_ (.A1(_1024_),
    .A2(\diff1_d[5] ),
    .B1(_1342_),
    .Y(_1347_));
 sky130_fd_sc_hd__a21oi_4 _4096_ (.A1(_1025_),
    .A2(\diff1_d[4] ),
    .B1(_1343_),
    .Y(_1348_));
 sky130_fd_sc_hd__nand2_1 _4097_ (.A(_1347_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__inv_2 _4098_ (.A(\diff1_d[3] ),
    .Y(_1350_));
 sky130_fd_sc_hd__nor2_1 _4099_ (.A(\diff1[3] ),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__a21oi_2 _4100_ (.A1(\diff1[3] ),
    .A2(_1350_),
    .B1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__inv_2 _4101_ (.A(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__a2bb2o_1 _4102_ (.A1_N(_1027_),
    .A2_N(\diff1_d[2] ),
    .B1(_1027_),
    .B2(\diff1_d[2] ),
    .X(_1354_));
 sky130_fd_sc_hd__inv_2 _4103_ (.A(\diff1_d[0] ),
    .Y(_1355_));
 sky130_fd_sc_hd__inv_2 _4104_ (.A(\diff1_d[1] ),
    .Y(_1356_));
 sky130_fd_sc_hd__o22a_1 _4105_ (.A1(_1030_),
    .A2(\diff1_d[1] ),
    .B1(\diff1[1] ),
    .B2(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__o21ai_1 _4106_ (.A1(\diff1[0] ),
    .A2(_1355_),
    .B1(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__o21ai_2 _4107_ (.A1(_1030_),
    .A2(\diff1_d[1] ),
    .B1(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__inv_2 _4108_ (.A(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__o32a_1 _4109_ (.A1(_1027_),
    .A2(\diff1_d[2] ),
    .A3(_1351_),
    .B1(_1026_),
    .B2(\diff1_d[3] ),
    .X(_1361_));
 sky130_fd_sc_hd__o31a_1 _4110_ (.A1(_1353_),
    .A2(_1354_),
    .A3(_1360_),
    .B1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__or4_4 _4111_ (.A(_1340_),
    .B(_1341_),
    .C(_1349_),
    .D(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__o311a_2 _4112_ (.A1(_1340_),
    .A2(_1341_),
    .A3(_1345_),
    .B1(_1346_),
    .C1(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__o22ai_1 _4113_ (.A1(_1014_),
    .A2(\diff1_d[13] ),
    .B1(_1015_),
    .B2(\diff1_d[12] ),
    .Y(_1365_));
 sky130_fd_sc_hd__o21ai_1 _4114_ (.A1(\diff1[13] ),
    .A2(_1322_),
    .B1(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__o22ai_1 _4115_ (.A1(_1019_),
    .A2(\diff1_d[9] ),
    .B1(_1020_),
    .B2(\diff1_d[8] ),
    .Y(_1367_));
 sky130_fd_sc_hd__o21ai_1 _4116_ (.A1(\diff1[9] ),
    .A2(_1331_),
    .B1(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__a211o_1 _4117_ (.A1(_1017_),
    .A2(\diff1_d[11] ),
    .B1(_1018_),
    .C1(\diff1_d[10] ),
    .X(_1369_));
 sky130_fd_sc_hd__o221a_1 _4118_ (.A1(_1017_),
    .A2(\diff1_d[11] ),
    .B1(_1330_),
    .B2(_1368_),
    .C1(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__o32a_1 _4119_ (.A1(_1013_),
    .A2(\diff1_d[14] ),
    .A3(_1317_),
    .B1(_1012_),
    .B2(\diff1_d[15] ),
    .X(_1371_));
 sky130_fd_sc_hd__o221a_1 _4120_ (.A1(_1321_),
    .A2(_1366_),
    .B1(_1327_),
    .B2(_1370_),
    .C1(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__o31a_2 _4121_ (.A1(_1327_),
    .A2(_1336_),
    .A3(_1364_),
    .B1(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__o22a_1 _4122_ (.A1(\diff1[17] ),
    .A2(_1305_),
    .B1(_1009_),
    .B2(\diff1_d[17] ),
    .X(_1374_));
 sky130_fd_sc_hd__inv_2 _4123_ (.A(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__o22a_1 _4124_ (.A1(_1011_),
    .A2(\diff1_d[16] ),
    .B1(\diff1[16] ),
    .B2(_1306_),
    .X(_1376_));
 sky130_fd_sc_hd__inv_2 _4125_ (.A(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__or2_1 _4126_ (.A(_1375_),
    .B(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__or2_1 _4127_ (.A(_1304_),
    .B(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__a21oi_2 _4128_ (.A1(\diff1[23] ),
    .A2(_1294_),
    .B1(_1295_),
    .Y(_1380_));
 sky130_fd_sc_hd__inv_2 _4129_ (.A(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__o2bb2a_1 _4130_ (.A1_N(_1003_),
    .A2_N(\diff1_d[22] ),
    .B1(_1002_),
    .B2(\diff1_d[22] ),
    .X(_1382_));
 sky130_fd_sc_hd__or4b_4 _4131_ (.A(_1379_),
    .B(_1381_),
    .C(_1300_),
    .D_N(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__o22a_2 _4132_ (.A1(_1295_),
    .A2(_1315_),
    .B1(_1373_),
    .B2(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__a2bb2o_1 _4133_ (.A1_N(_0994_),
    .A2_N(\diff1_d[28] ),
    .B1(\diff1[29] ),
    .B2(_1274_),
    .X(_1385_));
 sky130_fd_sc_hd__o21ai_1 _4134_ (.A1(\diff1[29] ),
    .A2(_1274_),
    .B1(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__o22ai_1 _4135_ (.A1(_0999_),
    .A2(\diff1_d[25] ),
    .B1(_1000_),
    .B2(\diff1_d[24] ),
    .Y(_1387_));
 sky130_fd_sc_hd__o21ai_1 _4136_ (.A1(\diff1[25] ),
    .A2(_1288_),
    .B1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__a211o_1 _4137_ (.A1(_0995_),
    .A2(\diff1_d[27] ),
    .B1(_0998_),
    .C1(\diff1_d[26] ),
    .X(_1389_));
 sky130_fd_sc_hd__o221a_1 _4138_ (.A1(_0995_),
    .A2(\diff1_d[27] ),
    .B1(_1287_),
    .B2(_1388_),
    .C1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__o32a_1 _4139_ (.A1(_0992_),
    .A2(\diff1_d[30] ),
    .A3(_1280_),
    .B1(_0991_),
    .B2(\diff1_d[31] ),
    .X(_1391_));
 sky130_fd_sc_hd__o221a_1 _4140_ (.A1(_1283_),
    .A2(_1386_),
    .B1(_1284_),
    .B2(_1390_),
    .C1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__o31a_1 _4141_ (.A1(_1284_),
    .A2(_1293_),
    .A3(_1384_),
    .B1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__o32a_1 _4142_ (.A1(_0989_),
    .A2(\diff1_d[32] ),
    .A3(_1269_),
    .B1(_0988_),
    .B2(\diff1_d[33] ),
    .X(_1394_));
 sky130_fd_sc_hd__o31a_1 _4143_ (.A1(_1271_),
    .A2(_1272_),
    .A3(_1393_),
    .B1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__o32a_1 _4144_ (.A1(_0987_),
    .A2(\diff1_d[34] ),
    .A3(_1264_),
    .B1(_0986_),
    .B2(\diff1_d[35] ),
    .X(_1396_));
 sky130_fd_sc_hd__o31a_1 _4145_ (.A1(_1266_),
    .A2(_1267_),
    .A3(_1395_),
    .B1(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__inv_2 _4146_ (.A(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__o221a_1 _4147_ (.A1(_1262_),
    .A2(_1397_),
    .B1(_1261_),
    .B2(_1398_),
    .C1(_1240_),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _4148_ (.A(_1395_),
    .B(_1267_),
    .X(_1399_));
 sky130_fd_sc_hd__o21ai_1 _4149_ (.A1(_0987_),
    .A2(\diff1_d[34] ),
    .B1(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__inv_2 _4150_ (.A(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__clkbuf_2 _4151_ (.A(_1239_),
    .X(_1402_));
 sky130_fd_sc_hd__o221a_1 _4152_ (.A1(_1266_),
    .A2(_1401_),
    .B1(_1265_),
    .B2(_1400_),
    .C1(_1402_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_2 _4153_ (.A(_0681_),
    .X(_1403_));
 sky130_fd_sc_hd__nand2_1 _4154_ (.A(_1395_),
    .B(_1267_),
    .Y(_1404_));
 sky130_fd_sc_hd__and3_1 _4155_ (.A(_1403_),
    .B(_1399_),
    .C(_1404_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _4156_ (.A(_1393_),
    .B(_1272_),
    .X(_1405_));
 sky130_fd_sc_hd__o21ai_1 _4157_ (.A1(_0989_),
    .A2(\diff1_d[32] ),
    .B1(_1405_),
    .Y(_1406_));
 sky130_fd_sc_hd__inv_2 _4158_ (.A(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__o221a_1 _4159_ (.A1(_1271_),
    .A2(_1407_),
    .B1(_1270_),
    .B2(_1406_),
    .C1(_1402_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2_1 _4160_ (.A(_1393_),
    .B(_1272_),
    .Y(_1408_));
 sky130_fd_sc_hd__and3_1 _4161_ (.A(_1403_),
    .B(_1405_),
    .C(_1408_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _4162_ (.A(_1278_),
    .Y(_1409_));
 sky130_fd_sc_hd__o21ai_1 _4163_ (.A1(_1384_),
    .A2(_1293_),
    .B1(_1390_),
    .Y(_1410_));
 sky130_fd_sc_hd__inv_2 _4164_ (.A(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__o21ai_1 _4165_ (.A1(_1277_),
    .A2(_1411_),
    .B1(_1386_),
    .Y(_1412_));
 sky130_fd_sc_hd__nand2_1 _4166_ (.A(_1409_),
    .B(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__o21ai_1 _4167_ (.A1(_0992_),
    .A2(\diff1_d[30] ),
    .B1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__inv_2 _4168_ (.A(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__o221a_1 _4169_ (.A1(_1282_),
    .A2(_1415_),
    .B1(_1281_),
    .B2(_1414_),
    .C1(_1402_),
    .X(_0290_));
 sky130_fd_sc_hd__o211a_1 _4170_ (.A1(_1409_),
    .A2(_1412_),
    .B1(_1241_),
    .C1(_1413_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _4171_ (.A(_1273_),
    .B(_1411_),
    .X(_1416_));
 sky130_fd_sc_hd__o21ai_1 _4172_ (.A1(_0994_),
    .A2(\diff1_d[28] ),
    .B1(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__inv_2 _4173_ (.A(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__o221a_1 _4174_ (.A1(_1276_),
    .A2(_1418_),
    .B1(_1275_),
    .B2(_1417_),
    .C1(_1402_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _4175_ (.A(_1273_),
    .Y(_1419_));
 sky130_fd_sc_hd__clkbuf_2 _4176_ (.A(_0679_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_2 _4177_ (.A(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__o211a_1 _4178_ (.A1(_1419_),
    .A2(_1410_),
    .B1(_1421_),
    .C1(_1416_),
    .X(_0287_));
 sky130_fd_sc_hd__inv_2 _4179_ (.A(_1286_),
    .Y(_1422_));
 sky130_fd_sc_hd__o21ai_1 _4180_ (.A1(_1384_),
    .A2(_1292_),
    .B1(_1388_),
    .Y(_1423_));
 sky130_fd_sc_hd__nand2_1 _4181_ (.A(_1422_),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__o21ai_1 _4182_ (.A1(_0998_),
    .A2(\diff1_d[26] ),
    .B1(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__inv_2 _4183_ (.A(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__inv_2 _4184_ (.A(_1285_),
    .Y(_1427_));
 sky130_fd_sc_hd__o221a_1 _4185_ (.A1(_1285_),
    .A2(_1426_),
    .B1(_1427_),
    .B2(_1425_),
    .C1(_1402_),
    .X(_0286_));
 sky130_fd_sc_hd__o211a_1 _4186_ (.A1(_1422_),
    .A2(_1423_),
    .B1(_1421_),
    .C1(_1424_),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _4187_ (.A(_1384_),
    .B(_1291_),
    .X(_1428_));
 sky130_fd_sc_hd__o21ai_1 _4188_ (.A1(_1000_),
    .A2(\diff1_d[24] ),
    .B1(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__inv_2 _4189_ (.A(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__buf_2 _4190_ (.A(_1239_),
    .X(_1431_));
 sky130_fd_sc_hd__o221a_1 _4191_ (.A1(_1290_),
    .A2(_1430_),
    .B1(_1289_),
    .B2(_1429_),
    .C1(_1431_),
    .X(_0284_));
 sky130_fd_sc_hd__nand2_1 _4192_ (.A(_1384_),
    .B(_1291_),
    .Y(_1432_));
 sky130_fd_sc_hd__and3_1 _4193_ (.A(_1403_),
    .B(_1428_),
    .C(_1432_),
    .X(_0283_));
 sky130_fd_sc_hd__o21ai_1 _4194_ (.A1(_1373_),
    .A2(_1379_),
    .B1(_1310_),
    .Y(_1433_));
 sky130_fd_sc_hd__inv_2 _4195_ (.A(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__o21ai_1 _4196_ (.A1(_1300_),
    .A2(_1434_),
    .B1(_1313_),
    .Y(_1435_));
 sky130_fd_sc_hd__nand2_1 _4197_ (.A(_1382_),
    .B(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hd__o21ai_1 _4198_ (.A1(_1003_),
    .A2(\diff1_d[22] ),
    .B1(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__inv_2 _4199_ (.A(_1437_),
    .Y(_1438_));
 sky130_fd_sc_hd__o221a_1 _4200_ (.A1(_1381_),
    .A2(_1438_),
    .B1(_1380_),
    .B2(_1437_),
    .C1(_1431_),
    .X(_0282_));
 sky130_fd_sc_hd__o211a_1 _4201_ (.A1(_1382_),
    .A2(_1435_),
    .B1(_1421_),
    .C1(_1436_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _4202_ (.A(_1299_),
    .B(_1434_),
    .X(_1439_));
 sky130_fd_sc_hd__o21ai_1 _4203_ (.A1(_1006_),
    .A2(\diff1_d[20] ),
    .B1(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__inv_2 _4204_ (.A(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__o221a_1 _4205_ (.A1(_1298_),
    .A2(_1441_),
    .B1(_1297_),
    .B2(_1440_),
    .C1(_1431_),
    .X(_0280_));
 sky130_fd_sc_hd__inv_2 _4206_ (.A(_1299_),
    .Y(_1442_));
 sky130_fd_sc_hd__o211a_1 _4207_ (.A1(_1442_),
    .A2(_1433_),
    .B1(_1421_),
    .C1(_1439_),
    .X(_0279_));
 sky130_fd_sc_hd__inv_2 _4208_ (.A(_1303_),
    .Y(_1443_));
 sky130_fd_sc_hd__o21ai_1 _4209_ (.A1(_1373_),
    .A2(_1378_),
    .B1(_1308_),
    .Y(_1444_));
 sky130_fd_sc_hd__nand2_1 _4210_ (.A(_1443_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__o21ai_1 _4211_ (.A1(_1008_),
    .A2(\diff1_d[18] ),
    .B1(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__inv_2 _4212_ (.A(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__o221a_1 _4213_ (.A1(_1302_),
    .A2(_1447_),
    .B1(_1301_),
    .B2(_1446_),
    .C1(_1431_),
    .X(_0278_));
 sky130_fd_sc_hd__o211a_1 _4214_ (.A1(_1443_),
    .A2(_1444_),
    .B1(_1421_),
    .C1(_1445_),
    .X(_0277_));
 sky130_fd_sc_hd__or2_1 _4215_ (.A(_1373_),
    .B(_1377_),
    .X(_1448_));
 sky130_fd_sc_hd__o21ai_1 _4216_ (.A1(_1011_),
    .A2(\diff1_d[16] ),
    .B1(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__inv_2 _4217_ (.A(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__o221a_1 _4218_ (.A1(_1375_),
    .A2(_1450_),
    .B1(_1374_),
    .B2(_1449_),
    .C1(_1431_),
    .X(_0276_));
 sky130_fd_sc_hd__inv_2 _4219_ (.A(_1373_),
    .Y(_1451_));
 sky130_fd_sc_hd__clkbuf_2 _4220_ (.A(_1420_),
    .X(_1452_));
 sky130_fd_sc_hd__o211a_1 _4221_ (.A1(_1451_),
    .A2(_1376_),
    .B1(_1452_),
    .C1(_1448_),
    .X(_0275_));
 sky130_fd_sc_hd__inv_2 _4222_ (.A(_1320_),
    .Y(_1453_));
 sky130_fd_sc_hd__o21ai_1 _4223_ (.A1(_1364_),
    .A2(_1336_),
    .B1(_1370_),
    .Y(_1454_));
 sky130_fd_sc_hd__inv_2 _4224_ (.A(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__o21ai_1 _4225_ (.A1(_1326_),
    .A2(_1455_),
    .B1(_1366_),
    .Y(_1456_));
 sky130_fd_sc_hd__nand2_1 _4226_ (.A(_1453_),
    .B(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__o21ai_1 _4227_ (.A1(_1013_),
    .A2(\diff1_d[14] ),
    .B1(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__inv_2 _4228_ (.A(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__clkbuf_2 _4229_ (.A(_1239_),
    .X(_1460_));
 sky130_fd_sc_hd__o221a_1 _4230_ (.A1(_1319_),
    .A2(_1459_),
    .B1(_1318_),
    .B2(_1458_),
    .C1(_1460_),
    .X(_0274_));
 sky130_fd_sc_hd__o211a_1 _4231_ (.A1(_1453_),
    .A2(_1456_),
    .B1(_1452_),
    .C1(_1457_),
    .X(_0273_));
 sky130_fd_sc_hd__or2_1 _4232_ (.A(_1325_),
    .B(_1455_),
    .X(_1461_));
 sky130_fd_sc_hd__o21ai_1 _4233_ (.A1(_1015_),
    .A2(\diff1_d[12] ),
    .B1(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__inv_2 _4234_ (.A(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__o221a_1 _4235_ (.A1(_1324_),
    .A2(_1463_),
    .B1(_1323_),
    .B2(_1462_),
    .C1(_1460_),
    .X(_0272_));
 sky130_fd_sc_hd__inv_2 _4236_ (.A(_1325_),
    .Y(_1464_));
 sky130_fd_sc_hd__o211a_1 _4237_ (.A1(_1464_),
    .A2(_1454_),
    .B1(_1452_),
    .C1(_1461_),
    .X(_0271_));
 sky130_fd_sc_hd__inv_2 _4238_ (.A(_1329_),
    .Y(_1465_));
 sky130_fd_sc_hd__o21ai_1 _4239_ (.A1(_1364_),
    .A2(_1335_),
    .B1(_1368_),
    .Y(_1466_));
 sky130_fd_sc_hd__nand2_1 _4240_ (.A(_1465_),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__o21ai_1 _4241_ (.A1(_1018_),
    .A2(\diff1_d[10] ),
    .B1(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__inv_2 _4242_ (.A(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _4243_ (.A(_1328_),
    .Y(_1470_));
 sky130_fd_sc_hd__o221a_1 _4244_ (.A1(_1328_),
    .A2(_1469_),
    .B1(_1470_),
    .B2(_1468_),
    .C1(_1460_),
    .X(_0270_));
 sky130_fd_sc_hd__o211a_1 _4245_ (.A1(_1465_),
    .A2(_1466_),
    .B1(_1452_),
    .C1(_1467_),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _4246_ (.A(_1364_),
    .B(_1334_),
    .X(_1471_));
 sky130_fd_sc_hd__o21ai_1 _4247_ (.A1(_1020_),
    .A2(\diff1_d[8] ),
    .B1(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__inv_2 _4248_ (.A(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__o221a_1 _4249_ (.A1(_1333_),
    .A2(_1473_),
    .B1(_1332_),
    .B2(_1472_),
    .C1(_1460_),
    .X(_0268_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(_1364_),
    .B(_1334_),
    .Y(_1474_));
 sky130_fd_sc_hd__and3_1 _4251_ (.A(_1403_),
    .B(_1471_),
    .C(_1474_),
    .X(_0267_));
 sky130_fd_sc_hd__inv_2 _4252_ (.A(_1341_),
    .Y(_1475_));
 sky130_fd_sc_hd__inv_2 _4253_ (.A(_1362_),
    .Y(_1476_));
 sky130_fd_sc_hd__a31o_1 _4254_ (.A1(_1347_),
    .A2(_1348_),
    .A3(_1476_),
    .B1(_1344_),
    .X(_1477_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(_1475_),
    .B(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__o21ai_1 _4256_ (.A1(_1023_),
    .A2(\diff1_d[6] ),
    .B1(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__inv_2 _4257_ (.A(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__o221a_1 _4258_ (.A1(_1340_),
    .A2(_1480_),
    .B1(_1339_),
    .B2(_1479_),
    .C1(_1460_),
    .X(_0266_));
 sky130_fd_sc_hd__o211a_1 _4259_ (.A1(_1475_),
    .A2(_1477_),
    .B1(_1452_),
    .C1(_1478_),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _4260_ (.A(_1476_),
    .B(_1348_),
    .Y(_1481_));
 sky130_fd_sc_hd__inv_2 _4261_ (.A(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__o21ai_1 _4262_ (.A1(_1343_),
    .A2(_1482_),
    .B1(_1347_),
    .Y(_1483_));
 sky130_fd_sc_hd__o311a_1 _4263_ (.A1(_1343_),
    .A2(_1482_),
    .A3(_1347_),
    .B1(_1254_),
    .C1(_1483_),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_4 _4264_ (.A(_1420_),
    .X(_1484_));
 sky130_fd_sc_hd__o211a_1 _4265_ (.A1(_1476_),
    .A2(_1348_),
    .B1(_1484_),
    .C1(_1481_),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _4266_ (.A(_1360_),
    .B(_1354_),
    .X(_1485_));
 sky130_fd_sc_hd__o21ai_1 _4267_ (.A1(_1027_),
    .A2(\diff1_d[2] ),
    .B1(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__inv_2 _4268_ (.A(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__clkbuf_4 _4269_ (.A(_1239_),
    .X(_1488_));
 sky130_fd_sc_hd__o221a_1 _4270_ (.A1(_1353_),
    .A2(_1487_),
    .B1(_1352_),
    .B2(_1486_),
    .C1(_1488_),
    .X(_0262_));
 sky130_fd_sc_hd__inv_2 _4271_ (.A(_1354_),
    .Y(_1489_));
 sky130_fd_sc_hd__o211a_1 _4272_ (.A1(_1359_),
    .A2(_1489_),
    .B1(_1484_),
    .C1(_1485_),
    .X(_0261_));
 sky130_fd_sc_hd__o311a_1 _4273_ (.A1(\diff1[0] ),
    .A2(_1355_),
    .A3(_1357_),
    .B1(_1254_),
    .C1(_1358_),
    .X(_0260_));
 sky130_fd_sc_hd__o22a_1 _4274_ (.A1(\diff1[0] ),
    .A2(_1355_),
    .B1(_1031_),
    .B2(\diff1_d[0] ),
    .X(_1490_));
 sky130_fd_sc_hd__nor2_1 _4275_ (.A(_1029_),
    .B(_1490_),
    .Y(_0259_));
 sky130_fd_sc_hd__a2bb2o_1 _4276_ (.A1_N(\acc3[36] ),
    .A2_N(\acc3_d2[36] ),
    .B1(\acc3[36] ),
    .B2(\acc3_d2[36] ),
    .X(_1491_));
 sky130_fd_sc_hd__inv_2 _4277_ (.A(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__inv_2 _4278_ (.A(\acc3_d2[35] ),
    .Y(_1493_));
 sky130_fd_sc_hd__nor2_1 _4279_ (.A(\acc3[35] ),
    .B(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__a21oi_2 _4280_ (.A1(\acc3[35] ),
    .A2(_1493_),
    .B1(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__inv_2 _4281_ (.A(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__inv_2 _4282_ (.A(\acc3[34] ),
    .Y(_1497_));
 sky130_fd_sc_hd__a2bb2o_1 _4283_ (.A1_N(_1497_),
    .A2_N(\acc3_d2[34] ),
    .B1(_1497_),
    .B2(\acc3_d2[34] ),
    .X(_1498_));
 sky130_fd_sc_hd__inv_2 _4284_ (.A(\acc3_d2[33] ),
    .Y(_1499_));
 sky130_fd_sc_hd__nor2_1 _4285_ (.A(\acc3[33] ),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__a21oi_2 _4286_ (.A1(\acc3[33] ),
    .A2(_1499_),
    .B1(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__inv_2 _4287_ (.A(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__inv_2 _4288_ (.A(\acc3[32] ),
    .Y(_1503_));
 sky130_fd_sc_hd__a2bb2o_1 _4289_ (.A1_N(_1503_),
    .A2_N(\acc3_d2[32] ),
    .B1(_1503_),
    .B2(\acc3_d2[32] ),
    .X(_1504_));
 sky130_fd_sc_hd__inv_2 _4290_ (.A(\acc3[28] ),
    .Y(_1505_));
 sky130_fd_sc_hd__buf_1 _4291_ (.A(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__a2bb2o_1 _4292_ (.A1_N(_1506_),
    .A2_N(\acc3_d2[28] ),
    .B1(_1505_),
    .B2(\acc3_d2[28] ),
    .X(_1507_));
 sky130_fd_sc_hd__inv_2 _4293_ (.A(\acc3[29] ),
    .Y(_1508_));
 sky130_fd_sc_hd__inv_2 _4294_ (.A(\acc3_d2[29] ),
    .Y(_1509_));
 sky130_fd_sc_hd__o22a_1 _4295_ (.A1(_1508_),
    .A2(\acc3_d2[29] ),
    .B1(\acc3[29] ),
    .B2(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__inv_2 _4296_ (.A(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__or2_1 _4297_ (.A(_1507_),
    .B(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__inv_2 _4298_ (.A(\acc3[30] ),
    .Y(_1513_));
 sky130_fd_sc_hd__a2bb2o_1 _4299_ (.A1_N(_1513_),
    .A2_N(\acc3_d2[30] ),
    .B1(_1513_),
    .B2(\acc3_d2[30] ),
    .X(_1514_));
 sky130_fd_sc_hd__inv_2 _4300_ (.A(\acc3_d2[31] ),
    .Y(_1515_));
 sky130_fd_sc_hd__nor2_1 _4301_ (.A(\acc3[31] ),
    .B(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__a21oi_2 _4302_ (.A1(\acc3[31] ),
    .A2(_1515_),
    .B1(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__inv_2 _4303_ (.A(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__or2_1 _4304_ (.A(_1514_),
    .B(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__or2_1 _4305_ (.A(_1512_),
    .B(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__inv_2 _4306_ (.A(\acc3[27] ),
    .Y(_1521_));
 sky130_fd_sc_hd__a2bb2o_1 _4307_ (.A1_N(_1521_),
    .A2_N(\acc3_d2[27] ),
    .B1(_1521_),
    .B2(\acc3_d2[27] ),
    .X(_1522_));
 sky130_fd_sc_hd__inv_2 _4308_ (.A(\acc3[26] ),
    .Y(_1523_));
 sky130_fd_sc_hd__a2bb2o_1 _4309_ (.A1_N(_1523_),
    .A2_N(\acc3_d2[26] ),
    .B1(_1523_),
    .B2(\acc3_d2[26] ),
    .X(_1524_));
 sky130_fd_sc_hd__or2_1 _4310_ (.A(_1522_),
    .B(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__inv_2 _4311_ (.A(\acc3[25] ),
    .Y(_1526_));
 sky130_fd_sc_hd__clkbuf_2 _4312_ (.A(\acc3[25] ),
    .X(_1527_));
 sky130_fd_sc_hd__inv_2 _4313_ (.A(\acc3_d2[25] ),
    .Y(_1528_));
 sky130_fd_sc_hd__o22a_1 _4314_ (.A1(_1526_),
    .A2(\acc3_d2[25] ),
    .B1(_1527_),
    .B2(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__inv_2 _4315_ (.A(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__inv_2 _4316_ (.A(\acc3[24] ),
    .Y(_1531_));
 sky130_fd_sc_hd__clkbuf_2 _4317_ (.A(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__a2bb2o_1 _4318_ (.A1_N(_1532_),
    .A2_N(\acc3_d2[24] ),
    .B1(_1531_),
    .B2(\acc3_d2[24] ),
    .X(_1533_));
 sky130_fd_sc_hd__or2_1 _4319_ (.A(_1530_),
    .B(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__or2_1 _4320_ (.A(_1525_),
    .B(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__inv_2 _4321_ (.A(\acc3_d2[23] ),
    .Y(_1536_));
 sky130_fd_sc_hd__nor2_1 _4322_ (.A(\acc3[23] ),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__inv_2 _4323_ (.A(\acc3[23] ),
    .Y(_1538_));
 sky130_fd_sc_hd__inv_2 _4324_ (.A(\acc3[22] ),
    .Y(_1539_));
 sky130_fd_sc_hd__buf_1 _4325_ (.A(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_2 _4326_ (.A(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_2 _4327_ (.A(\acc3[21] ),
    .X(_1542_));
 sky130_fd_sc_hd__inv_2 _4328_ (.A(\acc3_d2[21] ),
    .Y(_1543_));
 sky130_fd_sc_hd__inv_2 _4329_ (.A(\acc3[21] ),
    .Y(_1544_));
 sky130_fd_sc_hd__o22a_1 _4330_ (.A1(_1542_),
    .A2(_1543_),
    .B1(_1544_),
    .B2(\acc3_d2[21] ),
    .X(_1545_));
 sky130_fd_sc_hd__inv_2 _4331_ (.A(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__inv_2 _4332_ (.A(\acc3[20] ),
    .Y(_1547_));
 sky130_fd_sc_hd__buf_1 _4333_ (.A(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__a2bb2o_1 _4334_ (.A1_N(_1548_),
    .A2_N(\acc3_d2[20] ),
    .B1(_1547_),
    .B2(\acc3_d2[20] ),
    .X(_1549_));
 sky130_fd_sc_hd__or2_1 _4335_ (.A(_1546_),
    .B(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__inv_2 _4336_ (.A(\acc3[19] ),
    .Y(_1551_));
 sky130_fd_sc_hd__clkbuf_2 _4337_ (.A(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__o2bb2a_1 _4338_ (.A1_N(_1551_),
    .A2_N(\acc3_d2[19] ),
    .B1(_1551_),
    .B2(\acc3_d2[19] ),
    .X(_1553_));
 sky130_fd_sc_hd__inv_2 _4339_ (.A(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__inv_2 _4340_ (.A(\acc3[18] ),
    .Y(_1555_));
 sky130_fd_sc_hd__a2bb2o_1 _4341_ (.A1_N(_1555_),
    .A2_N(\acc3_d2[18] ),
    .B1(_1555_),
    .B2(\acc3_d2[18] ),
    .X(_1556_));
 sky130_fd_sc_hd__or2_1 _4342_ (.A(_1554_),
    .B(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_2 _4343_ (.A(\acc3[17] ),
    .X(_1558_));
 sky130_fd_sc_hd__inv_2 _4344_ (.A(\acc3_d2[17] ),
    .Y(_1559_));
 sky130_fd_sc_hd__inv_2 _4345_ (.A(\acc3_d2[16] ),
    .Y(_1560_));
 sky130_fd_sc_hd__a22o_1 _4346_ (.A1(\acc3[17] ),
    .A2(_1559_),
    .B1(\acc3[16] ),
    .B2(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__o21ai_1 _4347_ (.A1(_1558_),
    .A2(_1559_),
    .B1(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__clkbuf_2 _4348_ (.A(_1555_),
    .X(_1563_));
 sky130_fd_sc_hd__a211o_1 _4349_ (.A1(_1552_),
    .A2(\acc3_d2[19] ),
    .B1(_1563_),
    .C1(\acc3_d2[18] ),
    .X(_1564_));
 sky130_fd_sc_hd__o221a_1 _4350_ (.A1(_1552_),
    .A2(\acc3_d2[19] ),
    .B1(_1557_),
    .B2(_1562_),
    .C1(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__or2_1 _4351_ (.A(_1550_),
    .B(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__o22ai_1 _4352_ (.A1(_1544_),
    .A2(\acc3_d2[21] ),
    .B1(_1548_),
    .B2(\acc3_d2[20] ),
    .Y(_1567_));
 sky130_fd_sc_hd__o21ai_1 _4353_ (.A1(_1542_),
    .A2(_1543_),
    .B1(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__a22o_1 _4354_ (.A1(_1540_),
    .A2(\acc3_d2[22] ),
    .B1(_1566_),
    .B2(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__o221a_1 _4355_ (.A1(_1538_),
    .A2(\acc3_d2[23] ),
    .B1(_1541_),
    .B2(\acc3_d2[22] ),
    .C1(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__inv_2 _4356_ (.A(\acc3_d2[15] ),
    .Y(_1571_));
 sky130_fd_sc_hd__nor2_1 _4357_ (.A(\acc3[15] ),
    .B(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__a21oi_2 _4358_ (.A1(\acc3[15] ),
    .A2(_1571_),
    .B1(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__inv_2 _4359_ (.A(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__inv_2 _4360_ (.A(\acc3[14] ),
    .Y(_1575_));
 sky130_fd_sc_hd__a2bb2o_1 _4361_ (.A1_N(_1575_),
    .A2_N(\acc3_d2[14] ),
    .B1(_1575_),
    .B2(\acc3_d2[14] ),
    .X(_1576_));
 sky130_fd_sc_hd__or2_1 _4362_ (.A(_1574_),
    .B(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__inv_2 _4363_ (.A(\acc3[13] ),
    .Y(_1578_));
 sky130_fd_sc_hd__clkbuf_2 _4364_ (.A(\acc3[13] ),
    .X(_1579_));
 sky130_fd_sc_hd__inv_2 _4365_ (.A(\acc3_d2[13] ),
    .Y(_1580_));
 sky130_fd_sc_hd__o22a_1 _4366_ (.A1(_1578_),
    .A2(\acc3_d2[13] ),
    .B1(_1579_),
    .B2(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__inv_2 _4367_ (.A(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__inv_2 _4368_ (.A(\acc3[12] ),
    .Y(_1583_));
 sky130_fd_sc_hd__buf_1 _4369_ (.A(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__a2bb2o_1 _4370_ (.A1_N(_1584_),
    .A2_N(\acc3_d2[12] ),
    .B1(_1583_),
    .B2(\acc3_d2[12] ),
    .X(_1585_));
 sky130_fd_sc_hd__or2_1 _4371_ (.A(_1582_),
    .B(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__or2_1 _4372_ (.A(_1577_),
    .B(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__inv_2 _4373_ (.A(\acc3[11] ),
    .Y(_1588_));
 sky130_fd_sc_hd__a2bb2o_1 _4374_ (.A1_N(_1588_),
    .A2_N(\acc3_d2[11] ),
    .B1(_1588_),
    .B2(\acc3_d2[11] ),
    .X(_1589_));
 sky130_fd_sc_hd__inv_2 _4375_ (.A(\acc3[10] ),
    .Y(_1590_));
 sky130_fd_sc_hd__a2bb2o_1 _4376_ (.A1_N(_1590_),
    .A2_N(\acc3_d2[10] ),
    .B1(_1590_),
    .B2(\acc3_d2[10] ),
    .X(_1591_));
 sky130_fd_sc_hd__or2_1 _4377_ (.A(_1589_),
    .B(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__inv_2 _4378_ (.A(\acc3[9] ),
    .Y(_1593_));
 sky130_fd_sc_hd__clkbuf_2 _4379_ (.A(\acc3[9] ),
    .X(_1594_));
 sky130_fd_sc_hd__inv_2 _4380_ (.A(\acc3_d2[9] ),
    .Y(_1595_));
 sky130_fd_sc_hd__o22a_1 _4381_ (.A1(_1593_),
    .A2(\acc3_d2[9] ),
    .B1(_1594_),
    .B2(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__inv_2 _4382_ (.A(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(\acc3[8] ),
    .Y(_1598_));
 sky130_fd_sc_hd__buf_1 _4384_ (.A(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__a2bb2o_1 _4385_ (.A1_N(_1599_),
    .A2_N(\acc3_d2[8] ),
    .B1(_1598_),
    .B2(\acc3_d2[8] ),
    .X(_1600_));
 sky130_fd_sc_hd__or2_1 _4386_ (.A(_1597_),
    .B(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__or2_1 _4387_ (.A(_1592_),
    .B(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__inv_2 _4388_ (.A(\acc3_d2[7] ),
    .Y(_1603_));
 sky130_fd_sc_hd__nor2_1 _4389_ (.A(\acc3[7] ),
    .B(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__a21oi_2 _4390_ (.A1(\acc3[7] ),
    .A2(_1603_),
    .B1(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__inv_2 _4391_ (.A(_1605_),
    .Y(_1606_));
 sky130_fd_sc_hd__inv_2 _4392_ (.A(\acc3[6] ),
    .Y(_1607_));
 sky130_fd_sc_hd__a2bb2o_1 _4393_ (.A1_N(_1607_),
    .A2_N(\acc3_d2[6] ),
    .B1(_1607_),
    .B2(\acc3_d2[6] ),
    .X(_1608_));
 sky130_fd_sc_hd__inv_2 _4394_ (.A(\acc3[5] ),
    .Y(_1609_));
 sky130_fd_sc_hd__buf_2 _4395_ (.A(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__nor2_2 _4396_ (.A(_1609_),
    .B(\acc3_d2[5] ),
    .Y(_1611_));
 sky130_fd_sc_hd__clkinv_4 _4397_ (.A(\acc3[4] ),
    .Y(_1612_));
 sky130_fd_sc_hd__nor2_4 _4398_ (.A(_1612_),
    .B(\acc3_d2[4] ),
    .Y(_1613_));
 sky130_fd_sc_hd__o2bb2a_1 _4399_ (.A1_N(_1610_),
    .A2_N(\acc3_d2[5] ),
    .B1(_1611_),
    .B2(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__inv_2 _4400_ (.A(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__clkbuf_2 _4401_ (.A(_1607_),
    .X(_1616_));
 sky130_fd_sc_hd__inv_2 _4402_ (.A(\acc3[7] ),
    .Y(_1617_));
 sky130_fd_sc_hd__o32a_1 _4403_ (.A1(_1616_),
    .A2(\acc3_d2[6] ),
    .A3(_1604_),
    .B1(_1617_),
    .B2(\acc3_d2[7] ),
    .X(_1618_));
 sky130_fd_sc_hd__a21oi_4 _4404_ (.A1(_1610_),
    .A2(\acc3_d2[5] ),
    .B1(_1611_),
    .Y(_1619_));
 sky130_fd_sc_hd__a21oi_4 _4405_ (.A1(_1612_),
    .A2(\acc3_d2[4] ),
    .B1(_1613_),
    .Y(_1620_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_1619_),
    .B(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__inv_2 _4407_ (.A(\acc3_d2[3] ),
    .Y(_1622_));
 sky130_fd_sc_hd__nor2_1 _4408_ (.A(\acc3[3] ),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__a21oi_2 _4409_ (.A1(\acc3[3] ),
    .A2(_1622_),
    .B1(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__inv_2 _4410_ (.A(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__inv_2 _4411_ (.A(\acc3[2] ),
    .Y(_1626_));
 sky130_fd_sc_hd__a2bb2o_1 _4412_ (.A1_N(_1626_),
    .A2_N(\acc3_d2[2] ),
    .B1(_1626_),
    .B2(\acc3_d2[2] ),
    .X(_1627_));
 sky130_fd_sc_hd__inv_2 _4413_ (.A(\acc3[1] ),
    .Y(_1628_));
 sky130_fd_sc_hd__inv_2 _4414_ (.A(\acc3_d2[0] ),
    .Y(_1629_));
 sky130_fd_sc_hd__inv_2 _4415_ (.A(\acc3_d2[1] ),
    .Y(_1630_));
 sky130_fd_sc_hd__o22a_1 _4416_ (.A1(_1628_),
    .A2(\acc3_d2[1] ),
    .B1(\acc3[1] ),
    .B2(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__o21ai_1 _4417_ (.A1(\acc3[0] ),
    .A2(_1629_),
    .B1(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__o21ai_2 _4418_ (.A1(_1628_),
    .A2(\acc3_d2[1] ),
    .B1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__inv_2 _4419_ (.A(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4420_ (.A(_1626_),
    .X(_1635_));
 sky130_fd_sc_hd__inv_2 _4421_ (.A(\acc3[3] ),
    .Y(_1636_));
 sky130_fd_sc_hd__o32a_1 _4422_ (.A1(_1635_),
    .A2(\acc3_d2[2] ),
    .A3(_1623_),
    .B1(_1636_),
    .B2(\acc3_d2[3] ),
    .X(_1637_));
 sky130_fd_sc_hd__o31a_1 _4423_ (.A1(_1625_),
    .A2(_1627_),
    .A3(_1634_),
    .B1(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__or4_4 _4424_ (.A(_1606_),
    .B(_1608_),
    .C(_1621_),
    .D(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__o311a_2 _4425_ (.A1(_1606_),
    .A2(_1608_),
    .A3(_1615_),
    .B1(_1618_),
    .C1(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__o22ai_1 _4426_ (.A1(_1578_),
    .A2(\acc3_d2[13] ),
    .B1(_1584_),
    .B2(\acc3_d2[12] ),
    .Y(_1641_));
 sky130_fd_sc_hd__o21ai_1 _4427_ (.A1(_1579_),
    .A2(_1580_),
    .B1(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__clkbuf_2 _4428_ (.A(_1588_),
    .X(_1643_));
 sky130_fd_sc_hd__o22ai_1 _4429_ (.A1(_1593_),
    .A2(\acc3_d2[9] ),
    .B1(_1599_),
    .B2(\acc3_d2[8] ),
    .Y(_1644_));
 sky130_fd_sc_hd__o21ai_1 _4430_ (.A1(_1594_),
    .A2(_1595_),
    .B1(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__clkbuf_2 _4431_ (.A(_1590_),
    .X(_1646_));
 sky130_fd_sc_hd__a211o_1 _4432_ (.A1(_1643_),
    .A2(\acc3_d2[11] ),
    .B1(_1646_),
    .C1(\acc3_d2[10] ),
    .X(_1647_));
 sky130_fd_sc_hd__o221a_1 _4433_ (.A1(_1643_),
    .A2(\acc3_d2[11] ),
    .B1(_1592_),
    .B2(_1645_),
    .C1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_2 _4434_ (.A(_1575_),
    .X(_1649_));
 sky130_fd_sc_hd__inv_2 _4435_ (.A(\acc3[15] ),
    .Y(_1650_));
 sky130_fd_sc_hd__o32a_1 _4436_ (.A1(_1649_),
    .A2(\acc3_d2[14] ),
    .A3(_1572_),
    .B1(_1650_),
    .B2(\acc3_d2[15] ),
    .X(_1651_));
 sky130_fd_sc_hd__o221a_1 _4437_ (.A1(_1577_),
    .A2(_1642_),
    .B1(_1587_),
    .B2(_1648_),
    .C1(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__o31a_2 _4438_ (.A1(_1587_),
    .A2(_1602_),
    .A3(_1640_),
    .B1(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__inv_2 _4439_ (.A(\acc3[17] ),
    .Y(_1654_));
 sky130_fd_sc_hd__o22a_1 _4440_ (.A1(_1558_),
    .A2(_1559_),
    .B1(_1654_),
    .B2(\acc3_d2[17] ),
    .X(_1655_));
 sky130_fd_sc_hd__inv_2 _4441_ (.A(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__inv_2 _4442_ (.A(\acc3[16] ),
    .Y(_1657_));
 sky130_fd_sc_hd__o22a_1 _4443_ (.A1(_1657_),
    .A2(\acc3_d2[16] ),
    .B1(\acc3[16] ),
    .B2(_1560_),
    .X(_1658_));
 sky130_fd_sc_hd__inv_2 _4444_ (.A(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__or2_1 _4445_ (.A(_1656_),
    .B(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__or2_1 _4446_ (.A(_1557_),
    .B(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__a21oi_2 _4447_ (.A1(\acc3[23] ),
    .A2(_1536_),
    .B1(_1537_),
    .Y(_1662_));
 sky130_fd_sc_hd__inv_2 _4448_ (.A(_1662_),
    .Y(_1663_));
 sky130_fd_sc_hd__o2bb2a_1 _4449_ (.A1_N(_1540_),
    .A2_N(\acc3_d2[22] ),
    .B1(_1539_),
    .B2(\acc3_d2[22] ),
    .X(_1664_));
 sky130_fd_sc_hd__or4b_4 _4450_ (.A(_1661_),
    .B(_1663_),
    .C(_1550_),
    .D_N(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__o22a_2 _4451_ (.A1(_1537_),
    .A2(_1570_),
    .B1(_1653_),
    .B2(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_2 _4452_ (.A(\acc3[29] ),
    .X(_1667_));
 sky130_fd_sc_hd__a2bb2o_1 _4453_ (.A1_N(_1506_),
    .A2_N(\acc3_d2[28] ),
    .B1(_1667_),
    .B2(_1509_),
    .X(_1668_));
 sky130_fd_sc_hd__o21ai_1 _4454_ (.A1(_1667_),
    .A2(_1509_),
    .B1(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__clkbuf_2 _4455_ (.A(_1521_),
    .X(_1670_));
 sky130_fd_sc_hd__o22ai_1 _4456_ (.A1(_1526_),
    .A2(\acc3_d2[25] ),
    .B1(_1532_),
    .B2(\acc3_d2[24] ),
    .Y(_1671_));
 sky130_fd_sc_hd__o21ai_1 _4457_ (.A1(_1527_),
    .A2(_1528_),
    .B1(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__clkbuf_2 _4458_ (.A(_1523_),
    .X(_1673_));
 sky130_fd_sc_hd__a211o_1 _4459_ (.A1(_1670_),
    .A2(\acc3_d2[27] ),
    .B1(_1673_),
    .C1(\acc3_d2[26] ),
    .X(_1674_));
 sky130_fd_sc_hd__o221a_1 _4460_ (.A1(_1670_),
    .A2(\acc3_d2[27] ),
    .B1(_1525_),
    .B2(_1672_),
    .C1(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_2 _4461_ (.A(_1513_),
    .X(_1676_));
 sky130_fd_sc_hd__inv_2 _4462_ (.A(\acc3[31] ),
    .Y(_1677_));
 sky130_fd_sc_hd__o32a_1 _4463_ (.A1(_1676_),
    .A2(\acc3_d2[30] ),
    .A3(_1516_),
    .B1(_1677_),
    .B2(\acc3_d2[31] ),
    .X(_1678_));
 sky130_fd_sc_hd__o221a_1 _4464_ (.A1(_1519_),
    .A2(_1669_),
    .B1(_1520_),
    .B2(_1675_),
    .C1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__o31a_1 _4465_ (.A1(_1520_),
    .A2(_1535_),
    .A3(_1666_),
    .B1(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__clkbuf_2 _4466_ (.A(_1503_),
    .X(_1681_));
 sky130_fd_sc_hd__inv_2 _4467_ (.A(\acc3[33] ),
    .Y(_1682_));
 sky130_fd_sc_hd__o32a_1 _4468_ (.A1(_1681_),
    .A2(\acc3_d2[32] ),
    .A3(_1500_),
    .B1(_1682_),
    .B2(\acc3_d2[33] ),
    .X(_1683_));
 sky130_fd_sc_hd__o31a_1 _4469_ (.A1(_1502_),
    .A2(_1504_),
    .A3(_1680_),
    .B1(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_2 _4470_ (.A(_1497_),
    .X(_1685_));
 sky130_fd_sc_hd__inv_2 _4471_ (.A(\acc3[35] ),
    .Y(_1686_));
 sky130_fd_sc_hd__o32a_1 _4472_ (.A1(_1685_),
    .A2(\acc3_d2[34] ),
    .A3(_1494_),
    .B1(_1686_),
    .B2(\acc3_d2[35] ),
    .X(_1687_));
 sky130_fd_sc_hd__o31a_1 _4473_ (.A1(_1496_),
    .A2(_1498_),
    .A3(_1684_),
    .B1(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__inv_2 _4474_ (.A(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__o221a_1 _4475_ (.A1(_1492_),
    .A2(_1688_),
    .B1(_1491_),
    .B2(_1689_),
    .C1(_1488_),
    .X(_0258_));
 sky130_fd_sc_hd__or2_1 _4476_ (.A(_1684_),
    .B(_1498_),
    .X(_1690_));
 sky130_fd_sc_hd__o21ai_1 _4477_ (.A1(_1685_),
    .A2(\acc3_d2[34] ),
    .B1(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__inv_2 _4478_ (.A(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__o221a_1 _4479_ (.A1(_1496_),
    .A2(_1692_),
    .B1(_1495_),
    .B2(_1691_),
    .C1(_1488_),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(_1684_),
    .B(_1498_),
    .Y(_1693_));
 sky130_fd_sc_hd__and3_1 _4481_ (.A(_1403_),
    .B(_1690_),
    .C(_1693_),
    .X(_0256_));
 sky130_fd_sc_hd__or2_1 _4482_ (.A(_1680_),
    .B(_1504_),
    .X(_1694_));
 sky130_fd_sc_hd__o21ai_1 _4483_ (.A1(_1681_),
    .A2(\acc3_d2[32] ),
    .B1(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__inv_2 _4484_ (.A(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__o221a_1 _4485_ (.A1(_1502_),
    .A2(_1696_),
    .B1(_1501_),
    .B2(_1695_),
    .C1(_1488_),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _4486_ (.A(_1680_),
    .B(_1504_),
    .Y(_1697_));
 sky130_fd_sc_hd__and3_1 _4487_ (.A(_0767_),
    .B(_1694_),
    .C(_1697_),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _4488_ (.A(_1514_),
    .Y(_1698_));
 sky130_fd_sc_hd__o21ai_2 _4489_ (.A1(_1666_),
    .A2(_1535_),
    .B1(_1675_),
    .Y(_1699_));
 sky130_fd_sc_hd__inv_2 _4490_ (.A(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__o21ai_1 _4491_ (.A1(_1512_),
    .A2(_1700_),
    .B1(_1669_),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _4492_ (.A(_1698_),
    .B(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__o21ai_1 _4493_ (.A1(_1676_),
    .A2(\acc3_d2[30] ),
    .B1(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__inv_2 _4494_ (.A(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__o221a_1 _4495_ (.A1(_1518_),
    .A2(_1704_),
    .B1(_1517_),
    .B2(_1703_),
    .C1(_1488_),
    .X(_0253_));
 sky130_fd_sc_hd__o211a_1 _4496_ (.A1(_1698_),
    .A2(_1701_),
    .B1(_1484_),
    .C1(_1702_),
    .X(_0252_));
 sky130_fd_sc_hd__or2_1 _4497_ (.A(_1507_),
    .B(_1700_),
    .X(_1705_));
 sky130_fd_sc_hd__o21ai_1 _4498_ (.A1(_1506_),
    .A2(\acc3_d2[28] ),
    .B1(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__inv_2 _4499_ (.A(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__buf_1 _4500_ (.A(_0680_),
    .X(_1708_));
 sky130_fd_sc_hd__buf_2 _4501_ (.A(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__o221a_1 _4502_ (.A1(_1511_),
    .A2(_1707_),
    .B1(_1510_),
    .B2(_1706_),
    .C1(_1709_),
    .X(_0251_));
 sky130_fd_sc_hd__inv_2 _4503_ (.A(_1507_),
    .Y(_1710_));
 sky130_fd_sc_hd__o211a_1 _4504_ (.A1(_1710_),
    .A2(_1699_),
    .B1(_1484_),
    .C1(_1705_),
    .X(_0250_));
 sky130_fd_sc_hd__inv_2 _4505_ (.A(_1524_),
    .Y(_1711_));
 sky130_fd_sc_hd__o21ai_1 _4506_ (.A1(_1666_),
    .A2(_1534_),
    .B1(_1672_),
    .Y(_1712_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(_1711_),
    .B(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__o21ai_1 _4508_ (.A1(_1673_),
    .A2(\acc3_d2[26] ),
    .B1(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__inv_2 _4509_ (.A(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__inv_2 _4510_ (.A(_1522_),
    .Y(_1716_));
 sky130_fd_sc_hd__o221a_1 _4511_ (.A1(_1522_),
    .A2(_1715_),
    .B1(_1716_),
    .B2(_1714_),
    .C1(_1709_),
    .X(_0249_));
 sky130_fd_sc_hd__o211a_1 _4512_ (.A1(_1711_),
    .A2(_1712_),
    .B1(_1484_),
    .C1(_1713_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _4513_ (.A(_1666_),
    .B(_1533_),
    .X(_1717_));
 sky130_fd_sc_hd__o21ai_1 _4514_ (.A1(_1532_),
    .A2(\acc3_d2[24] ),
    .B1(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__inv_2 _4515_ (.A(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__o221a_1 _4516_ (.A1(_1530_),
    .A2(_1719_),
    .B1(_1529_),
    .B2(_1718_),
    .C1(_1709_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_1666_),
    .B(_1533_),
    .Y(_1720_));
 sky130_fd_sc_hd__and3_1 _4518_ (.A(_0767_),
    .B(_1717_),
    .C(_1720_),
    .X(_0246_));
 sky130_fd_sc_hd__o21ai_1 _4519_ (.A1(_1653_),
    .A2(_1661_),
    .B1(_1565_),
    .Y(_1721_));
 sky130_fd_sc_hd__inv_2 _4520_ (.A(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__o21ai_1 _4521_ (.A1(_1550_),
    .A2(_1722_),
    .B1(_1568_),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_1 _4522_ (.A(_1664_),
    .B(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__o21ai_1 _4523_ (.A1(_1541_),
    .A2(\acc3_d2[22] ),
    .B1(_1724_),
    .Y(_1725_));
 sky130_fd_sc_hd__inv_2 _4524_ (.A(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__o221a_1 _4525_ (.A1(_1663_),
    .A2(_1726_),
    .B1(_1662_),
    .B2(_1725_),
    .C1(_1709_),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_2 _4526_ (.A(_1420_),
    .X(_1727_));
 sky130_fd_sc_hd__o211a_1 _4527_ (.A1(_1664_),
    .A2(_1723_),
    .B1(_1727_),
    .C1(_1724_),
    .X(_0244_));
 sky130_fd_sc_hd__or2_1 _4528_ (.A(_1549_),
    .B(_1722_),
    .X(_1728_));
 sky130_fd_sc_hd__o21ai_1 _4529_ (.A1(_1548_),
    .A2(\acc3_d2[20] ),
    .B1(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hd__inv_2 _4530_ (.A(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__o221a_1 _4531_ (.A1(_1546_),
    .A2(_1730_),
    .B1(_1545_),
    .B2(_1729_),
    .C1(_1709_),
    .X(_0243_));
 sky130_fd_sc_hd__inv_2 _4532_ (.A(_1549_),
    .Y(_1731_));
 sky130_fd_sc_hd__o211a_1 _4533_ (.A1(_1731_),
    .A2(_1721_),
    .B1(_1727_),
    .C1(_1728_),
    .X(_0242_));
 sky130_fd_sc_hd__inv_2 _4534_ (.A(_1556_),
    .Y(_1732_));
 sky130_fd_sc_hd__o21ai_1 _4535_ (.A1(_1653_),
    .A2(_1660_),
    .B1(_1562_),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(_1732_),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__o21ai_1 _4537_ (.A1(_1563_),
    .A2(\acc3_d2[18] ),
    .B1(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__inv_2 _4538_ (.A(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__clkbuf_2 _4539_ (.A(_1708_),
    .X(_1737_));
 sky130_fd_sc_hd__o221a_1 _4540_ (.A1(_1554_),
    .A2(_1736_),
    .B1(_1553_),
    .B2(_1735_),
    .C1(_1737_),
    .X(_0241_));
 sky130_fd_sc_hd__o211a_1 _4541_ (.A1(_1732_),
    .A2(_1733_),
    .B1(_1727_),
    .C1(_1734_),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _4542_ (.A(_1653_),
    .B(_1659_),
    .X(_1738_));
 sky130_fd_sc_hd__o21ai_1 _4543_ (.A1(_1657_),
    .A2(\acc3_d2[16] ),
    .B1(_1738_),
    .Y(_1739_));
 sky130_fd_sc_hd__inv_2 _4544_ (.A(_1739_),
    .Y(_1740_));
 sky130_fd_sc_hd__o221a_1 _4545_ (.A1(_1656_),
    .A2(_1740_),
    .B1(_1655_),
    .B2(_1739_),
    .C1(_1737_),
    .X(_0239_));
 sky130_fd_sc_hd__inv_2 _4546_ (.A(_1653_),
    .Y(_1741_));
 sky130_fd_sc_hd__o211a_1 _4547_ (.A1(_1741_),
    .A2(_1658_),
    .B1(_1727_),
    .C1(_1738_),
    .X(_0238_));
 sky130_fd_sc_hd__inv_2 _4548_ (.A(_1576_),
    .Y(_1742_));
 sky130_fd_sc_hd__o21ai_1 _4549_ (.A1(_1640_),
    .A2(_1602_),
    .B1(_1648_),
    .Y(_1743_));
 sky130_fd_sc_hd__inv_2 _4550_ (.A(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__o21ai_1 _4551_ (.A1(_1586_),
    .A2(_1744_),
    .B1(_1642_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(_1742_),
    .B(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__o21ai_1 _4553_ (.A1(_1649_),
    .A2(\acc3_d2[14] ),
    .B1(_1746_),
    .Y(_1747_));
 sky130_fd_sc_hd__inv_2 _4554_ (.A(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__o221a_1 _4555_ (.A1(_1574_),
    .A2(_1748_),
    .B1(_1573_),
    .B2(_1747_),
    .C1(_1737_),
    .X(_0237_));
 sky130_fd_sc_hd__o211a_1 _4556_ (.A1(_1742_),
    .A2(_1745_),
    .B1(_1727_),
    .C1(_1746_),
    .X(_0236_));
 sky130_fd_sc_hd__or2_1 _4557_ (.A(_1585_),
    .B(_1744_),
    .X(_1749_));
 sky130_fd_sc_hd__o21ai_1 _4558_ (.A1(_1584_),
    .A2(\acc3_d2[12] ),
    .B1(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__inv_2 _4559_ (.A(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__o221a_1 _4560_ (.A1(_1582_),
    .A2(_1751_),
    .B1(_1581_),
    .B2(_1750_),
    .C1(_1737_),
    .X(_0235_));
 sky130_fd_sc_hd__inv_2 _4561_ (.A(_1585_),
    .Y(_1752_));
 sky130_fd_sc_hd__clkbuf_2 _4562_ (.A(_1420_),
    .X(_1753_));
 sky130_fd_sc_hd__o211a_1 _4563_ (.A1(_1752_),
    .A2(_1743_),
    .B1(_1753_),
    .C1(_1749_),
    .X(_0234_));
 sky130_fd_sc_hd__inv_2 _4564_ (.A(_1591_),
    .Y(_1754_));
 sky130_fd_sc_hd__o21ai_1 _4565_ (.A1(_1640_),
    .A2(_1601_),
    .B1(_1645_),
    .Y(_1755_));
 sky130_fd_sc_hd__nand2_1 _4566_ (.A(_1754_),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__o21ai_1 _4567_ (.A1(_1646_),
    .A2(\acc3_d2[10] ),
    .B1(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__inv_2 _4568_ (.A(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__inv_2 _4569_ (.A(_1589_),
    .Y(_1759_));
 sky130_fd_sc_hd__o221a_1 _4570_ (.A1(_1589_),
    .A2(_1758_),
    .B1(_1759_),
    .B2(_1757_),
    .C1(_1737_),
    .X(_0233_));
 sky130_fd_sc_hd__o211a_1 _4571_ (.A1(_1754_),
    .A2(_1755_),
    .B1(_1753_),
    .C1(_1756_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _4572_ (.A(_1640_),
    .B(_1600_),
    .X(_1760_));
 sky130_fd_sc_hd__o21ai_1 _4573_ (.A1(_1599_),
    .A2(\acc3_d2[8] ),
    .B1(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__inv_2 _4574_ (.A(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__buf_2 _4575_ (.A(_1708_),
    .X(_1763_));
 sky130_fd_sc_hd__o221a_1 _4576_ (.A1(_1597_),
    .A2(_1762_),
    .B1(_1596_),
    .B2(_1761_),
    .C1(_1763_),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_1640_),
    .B(_1600_),
    .Y(_1764_));
 sky130_fd_sc_hd__and3_1 _4578_ (.A(_0767_),
    .B(_1760_),
    .C(_1764_),
    .X(_0230_));
 sky130_fd_sc_hd__inv_2 _4579_ (.A(_1608_),
    .Y(_1765_));
 sky130_fd_sc_hd__inv_2 _4580_ (.A(_1638_),
    .Y(_1766_));
 sky130_fd_sc_hd__a31o_1 _4581_ (.A1(_1619_),
    .A2(_1620_),
    .A3(_1766_),
    .B1(_1614_),
    .X(_1767_));
 sky130_fd_sc_hd__nand2_1 _4582_ (.A(_1765_),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__o21ai_1 _4583_ (.A1(_1616_),
    .A2(\acc3_d2[6] ),
    .B1(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__inv_2 _4584_ (.A(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__o221a_1 _4585_ (.A1(_1606_),
    .A2(_1770_),
    .B1(_1605_),
    .B2(_1769_),
    .C1(_1763_),
    .X(_0229_));
 sky130_fd_sc_hd__o211a_1 _4586_ (.A1(_1765_),
    .A2(_1767_),
    .B1(_1753_),
    .C1(_1768_),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_1 _4587_ (.A(_1766_),
    .B(_1620_),
    .Y(_1771_));
 sky130_fd_sc_hd__inv_2 _4588_ (.A(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__o21ai_1 _4589_ (.A1(_1613_),
    .A2(_1772_),
    .B1(_1619_),
    .Y(_1773_));
 sky130_fd_sc_hd__o311a_1 _4590_ (.A1(_1613_),
    .A2(_1772_),
    .A3(_1619_),
    .B1(_1254_),
    .C1(_1773_),
    .X(_0227_));
 sky130_fd_sc_hd__o211a_1 _4591_ (.A1(_1766_),
    .A2(_1620_),
    .B1(_1753_),
    .C1(_1771_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _4592_ (.A(_1634_),
    .B(_1627_),
    .X(_1774_));
 sky130_fd_sc_hd__o21ai_1 _4593_ (.A1(_1635_),
    .A2(\acc3_d2[2] ),
    .B1(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__inv_2 _4594_ (.A(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__o221a_1 _4595_ (.A1(_1625_),
    .A2(_1776_),
    .B1(_1624_),
    .B2(_1775_),
    .C1(_1763_),
    .X(_0225_));
 sky130_fd_sc_hd__inv_2 _4596_ (.A(_1627_),
    .Y(_1777_));
 sky130_fd_sc_hd__o211a_1 _4597_ (.A1(_1633_),
    .A2(_1777_),
    .B1(_1753_),
    .C1(_1774_),
    .X(_0224_));
 sky130_fd_sc_hd__o311a_1 _4598_ (.A1(\acc3[0] ),
    .A2(_1629_),
    .A3(_1631_),
    .B1(_0688_),
    .C1(_1632_),
    .X(_0223_));
 sky130_fd_sc_hd__inv_2 _4599_ (.A(\acc3[0] ),
    .Y(_1778_));
 sky130_fd_sc_hd__o22a_1 _4600_ (.A1(\acc3[0] ),
    .A2(_1629_),
    .B1(_1778_),
    .B2(\acc3_d2[0] ),
    .X(_1779_));
 sky130_fd_sc_hd__nor2_1 _4601_ (.A(_1029_),
    .B(_1779_),
    .Y(_0222_));
 sky130_fd_sc_hd__clkbuf_2 _4602_ (.A(_1028_),
    .X(_1780_));
 sky130_fd_sc_hd__inv_2 _4603_ (.A(\acc3[36] ),
    .Y(_1781_));
 sky130_fd_sc_hd__nor2_1 _4604_ (.A(_1780_),
    .B(_1781_),
    .Y(_0221_));
 sky130_fd_sc_hd__nor2_1 _4605_ (.A(_1780_),
    .B(_1686_),
    .Y(_0220_));
 sky130_fd_sc_hd__nor2_1 _4606_ (.A(_1780_),
    .B(_1685_),
    .Y(_0219_));
 sky130_fd_sc_hd__nor2_1 _4607_ (.A(_1780_),
    .B(_1682_),
    .Y(_0218_));
 sky130_fd_sc_hd__nor2_1 _4608_ (.A(_1780_),
    .B(_1681_),
    .Y(_0217_));
 sky130_fd_sc_hd__clkbuf_2 _4609_ (.A(_1028_),
    .X(_1782_));
 sky130_fd_sc_hd__nor2_1 _4610_ (.A(_1782_),
    .B(_1677_),
    .Y(_0216_));
 sky130_fd_sc_hd__nor2_1 _4611_ (.A(_1782_),
    .B(_1676_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _4612_ (.A(_1782_),
    .B(_1508_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _4613_ (.A(_1782_),
    .B(_1506_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _4614_ (.A(_1782_),
    .B(_1670_),
    .Y(_0212_));
 sky130_fd_sc_hd__buf_2 _4615_ (.A(_1028_),
    .X(_1783_));
 sky130_fd_sc_hd__nor2_1 _4616_ (.A(_1783_),
    .B(_1673_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor2_1 _4617_ (.A(_1783_),
    .B(_1526_),
    .Y(_0210_));
 sky130_fd_sc_hd__nor2_1 _4618_ (.A(_1783_),
    .B(_1532_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _4619_ (.A(_1783_),
    .B(_1538_),
    .Y(_0208_));
 sky130_fd_sc_hd__nor2_1 _4620_ (.A(_1783_),
    .B(_1541_),
    .Y(_0207_));
 sky130_fd_sc_hd__clkbuf_2 _4621_ (.A(_1028_),
    .X(_1784_));
 sky130_fd_sc_hd__nor2_1 _4622_ (.A(_1784_),
    .B(_1544_),
    .Y(_0206_));
 sky130_fd_sc_hd__nor2_1 _4623_ (.A(_1784_),
    .B(_1548_),
    .Y(_0205_));
 sky130_fd_sc_hd__nor2_1 _4624_ (.A(_1784_),
    .B(_1552_),
    .Y(_0204_));
 sky130_fd_sc_hd__nor2_1 _4625_ (.A(_1784_),
    .B(_1563_),
    .Y(_0203_));
 sky130_fd_sc_hd__nor2_1 _4626_ (.A(_1784_),
    .B(_1654_),
    .Y(_0202_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4627_ (.A(_0817_),
    .X(_1785_));
 sky130_fd_sc_hd__nor2_1 _4628_ (.A(_1785_),
    .B(_1657_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor2_1 _4629_ (.A(_1785_),
    .B(_1650_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _4630_ (.A(_1785_),
    .B(_1649_),
    .Y(_0199_));
 sky130_fd_sc_hd__nor2_1 _4631_ (.A(_1785_),
    .B(_1578_),
    .Y(_0198_));
 sky130_fd_sc_hd__nor2_1 _4632_ (.A(_1785_),
    .B(_1584_),
    .Y(_0197_));
 sky130_fd_sc_hd__clkbuf_2 _4633_ (.A(_0817_),
    .X(_1786_));
 sky130_fd_sc_hd__nor2_1 _4634_ (.A(_1786_),
    .B(_1643_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _4635_ (.A(_1786_),
    .B(_1646_),
    .Y(_0195_));
 sky130_fd_sc_hd__nor2_1 _4636_ (.A(_1786_),
    .B(_1593_),
    .Y(_0194_));
 sky130_fd_sc_hd__nor2_1 _4637_ (.A(_1786_),
    .B(_1599_),
    .Y(_0193_));
 sky130_fd_sc_hd__nor2_1 _4638_ (.A(_1786_),
    .B(_1617_),
    .Y(_0192_));
 sky130_fd_sc_hd__clkbuf_2 _4639_ (.A(_0817_),
    .X(_1787_));
 sky130_fd_sc_hd__nor2_1 _4640_ (.A(_1787_),
    .B(_1616_),
    .Y(_0191_));
 sky130_fd_sc_hd__nor2_1 _4641_ (.A(_1787_),
    .B(_1610_),
    .Y(_0190_));
 sky130_fd_sc_hd__nor2_1 _4642_ (.A(_1787_),
    .B(_1612_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _4643_ (.A(_1787_),
    .B(_1636_),
    .Y(_0188_));
 sky130_fd_sc_hd__nor2_1 _4644_ (.A(_1787_),
    .B(_1635_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _4645_ (.A(_0814_),
    .B(_1628_),
    .Y(_0186_));
 sky130_fd_sc_hd__nor2_1 _4646_ (.A(_0814_),
    .B(_1778_),
    .Y(_0185_));
 sky130_fd_sc_hd__nor2_1 _4647_ (.A(_0814_),
    .B(_2323_),
    .Y(_0184_));
 sky130_fd_sc_hd__buf_1 _4648_ (.A(_0847_),
    .X(_0072_));
 sky130_fd_sc_hd__o22a_1 _4649_ (.A1(\acc3[36] ),
    .A2(\acc2[36] ),
    .B1(_1781_),
    .B2(_2328_),
    .X(_1788_));
 sky130_fd_sc_hd__nor2_1 _4650_ (.A(\acc3[35] ),
    .B(\acc2[35] ),
    .Y(_1789_));
 sky130_fd_sc_hd__a21oi_2 _4651_ (.A1(\acc3[35] ),
    .A2(\acc2[35] ),
    .B1(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__inv_2 _4652_ (.A(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__o22a_1 _4653_ (.A1(_1497_),
    .A2(_2334_),
    .B1(\acc3[34] ),
    .B2(\acc2[34] ),
    .X(_1792_));
 sky130_fd_sc_hd__inv_2 _4654_ (.A(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__nor2_1 _4655_ (.A(\acc3[33] ),
    .B(\acc2[33] ),
    .Y(_1794_));
 sky130_fd_sc_hd__a21oi_2 _4656_ (.A1(\acc3[33] ),
    .A2(\acc2[33] ),
    .B1(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__inv_2 _4657_ (.A(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__o22a_1 _4658_ (.A1(_1503_),
    .A2(_2342_),
    .B1(\acc3[32] ),
    .B2(\acc2[32] ),
    .X(_1797_));
 sky130_fd_sc_hd__inv_2 _4659_ (.A(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__o22a_1 _4660_ (.A1(\acc3[28] ),
    .A2(\acc2[28] ),
    .B1(_1505_),
    .B2(_2347_),
    .X(_1799_));
 sky130_fd_sc_hd__inv_2 _4661_ (.A(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__o22a_1 _4662_ (.A1(_1667_),
    .A2(\acc2[29] ),
    .B1(_1508_),
    .B2(_2352_),
    .X(_1801_));
 sky130_fd_sc_hd__inv_2 _4663_ (.A(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__or2_1 _4664_ (.A(_1800_),
    .B(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__o22a_1 _4665_ (.A1(\acc3[30] ),
    .A2(\acc2[30] ),
    .B1(_1513_),
    .B2(_2357_),
    .X(_1804_));
 sky130_fd_sc_hd__nor2_1 _4666_ (.A(\acc3[31] ),
    .B(\acc2[31] ),
    .Y(_1805_));
 sky130_fd_sc_hd__a21oi_2 _4667_ (.A1(\acc3[31] ),
    .A2(\acc2[31] ),
    .B1(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _4668_ (.A(_1804_),
    .B(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__or2_1 _4669_ (.A(_1803_),
    .B(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__o22a_1 _4670_ (.A1(_1521_),
    .A2(_2365_),
    .B1(\acc3[27] ),
    .B2(\acc2[27] ),
    .X(_1809_));
 sky130_fd_sc_hd__o22a_1 _4671_ (.A1(_1523_),
    .A2(_2369_),
    .B1(\acc3[26] ),
    .B2(\acc2[26] ),
    .X(_1810_));
 sky130_fd_sc_hd__nand2_1 _4672_ (.A(_1809_),
    .B(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__o22a_1 _4673_ (.A1(_1526_),
    .A2(_0503_),
    .B1(_1527_),
    .B2(\acc2[25] ),
    .X(_1812_));
 sky130_fd_sc_hd__inv_2 _4674_ (.A(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__o22a_1 _4675_ (.A1(_1531_),
    .A2(_0508_),
    .B1(\acc3[24] ),
    .B2(\acc2[24] ),
    .X(_1814_));
 sky130_fd_sc_hd__inv_2 _4676_ (.A(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__or2_1 _4677_ (.A(_1813_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__or2_1 _4678_ (.A(_1811_),
    .B(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__nor2_2 _4679_ (.A(\acc3[23] ),
    .B(\acc2[23] ),
    .Y(_1818_));
 sky130_fd_sc_hd__o22a_1 _4680_ (.A1(_1542_),
    .A2(\acc2[21] ),
    .B1(_1544_),
    .B2(_0521_),
    .X(_1819_));
 sky130_fd_sc_hd__inv_2 _4681_ (.A(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__o22a_1 _4682_ (.A1(_1547_),
    .A2(_0525_),
    .B1(\acc3[20] ),
    .B2(\acc2[20] ),
    .X(_1821_));
 sky130_fd_sc_hd__inv_2 _4683_ (.A(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__or2_1 _4684_ (.A(_1820_),
    .B(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__o22a_1 _4685_ (.A1(\acc3[19] ),
    .A2(\acc2[19] ),
    .B1(_1551_),
    .B2(_0530_),
    .X(_1824_));
 sky130_fd_sc_hd__o22a_1 _4686_ (.A1(_1555_),
    .A2(_0534_),
    .B1(\acc3[18] ),
    .B2(\acc2[18] ),
    .X(_1825_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_1824_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__a22o_1 _4688_ (.A1(_1558_),
    .A2(\acc2[17] ),
    .B1(\acc3[16] ),
    .B2(\acc2[16] ),
    .X(_1827_));
 sky130_fd_sc_hd__o21ai_1 _4689_ (.A1(_1558_),
    .A2(_0538_),
    .B1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__a211o_1 _4690_ (.A1(_1552_),
    .A2(_0531_),
    .B1(_1563_),
    .C1(_0535_),
    .X(_1829_));
 sky130_fd_sc_hd__o221a_1 _4691_ (.A1(_1552_),
    .A2(_0531_),
    .B1(_1826_),
    .B2(_1828_),
    .C1(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__or2_1 _4692_ (.A(_1823_),
    .B(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__a22o_1 _4693_ (.A1(_1542_),
    .A2(_0519_),
    .B1(\acc3[20] ),
    .B2(\acc2[20] ),
    .X(_1832_));
 sky130_fd_sc_hd__o21ai_1 _4694_ (.A1(_1542_),
    .A2(_0519_),
    .B1(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__a22o_1 _4695_ (.A1(_1540_),
    .A2(_0517_),
    .B1(_1831_),
    .B2(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__o221a_1 _4696_ (.A1(_1538_),
    .A2(_0515_),
    .B1(_1541_),
    .B2(_0518_),
    .C1(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__nor2_1 _4697_ (.A(\acc3[15] ),
    .B(\acc2[15] ),
    .Y(_1836_));
 sky130_fd_sc_hd__a21oi_2 _4698_ (.A1(\acc3[15] ),
    .A2(\acc2[15] ),
    .B1(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__o22a_1 _4699_ (.A1(_1575_),
    .A2(_0551_),
    .B1(\acc3[14] ),
    .B2(\acc2[14] ),
    .X(_1838_));
 sky130_fd_sc_hd__nand2_1 _4700_ (.A(_1837_),
    .B(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__o22a_1 _4701_ (.A1(_1578_),
    .A2(_0556_),
    .B1(_1579_),
    .B2(\acc2[13] ),
    .X(_1840_));
 sky130_fd_sc_hd__inv_2 _4702_ (.A(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__o22a_1 _4703_ (.A1(_1583_),
    .A2(_0561_),
    .B1(\acc3[12] ),
    .B2(\acc2[12] ),
    .X(_1842_));
 sky130_fd_sc_hd__inv_2 _4704_ (.A(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__or2_1 _4705_ (.A(_1841_),
    .B(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__or2_1 _4706_ (.A(_1839_),
    .B(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__o22a_1 _4707_ (.A1(_1588_),
    .A2(_0567_),
    .B1(\acc3[11] ),
    .B2(\acc2[11] ),
    .X(_1846_));
 sky130_fd_sc_hd__o22a_1 _4708_ (.A1(_1590_),
    .A2(_0571_),
    .B1(\acc3[10] ),
    .B2(\acc2[10] ),
    .X(_1847_));
 sky130_fd_sc_hd__nand2_1 _4709_ (.A(_1846_),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__o22a_1 _4710_ (.A1(_1593_),
    .A2(_0576_),
    .B1(_1594_),
    .B2(\acc2[9] ),
    .X(_1849_));
 sky130_fd_sc_hd__inv_2 _4711_ (.A(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__o22a_1 _4712_ (.A1(_1598_),
    .A2(_0581_),
    .B1(\acc3[8] ),
    .B2(\acc2[8] ),
    .X(_1851_));
 sky130_fd_sc_hd__inv_2 _4713_ (.A(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__or2_1 _4714_ (.A(_1850_),
    .B(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__or2_1 _4715_ (.A(_1848_),
    .B(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__nor2_1 _4716_ (.A(\acc3[7] ),
    .B(\acc2[7] ),
    .Y(_1855_));
 sky130_fd_sc_hd__a21oi_2 _4717_ (.A1(\acc3[7] ),
    .A2(\acc2[7] ),
    .B1(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__inv_2 _4718_ (.A(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__o22a_1 _4719_ (.A1(_1607_),
    .A2(_0590_),
    .B1(\acc3[6] ),
    .B2(\acc2[6] ),
    .X(_1858_));
 sky130_fd_sc_hd__inv_2 _4720_ (.A(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__nor2_2 _4721_ (.A(_1610_),
    .B(_0595_),
    .Y(_1860_));
 sky130_fd_sc_hd__nor2_4 _4722_ (.A(_1612_),
    .B(_0598_),
    .Y(_1861_));
 sky130_fd_sc_hd__o22a_1 _4723_ (.A1(\acc3[5] ),
    .A2(\acc2[5] ),
    .B1(_1860_),
    .B2(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__inv_2 _4724_ (.A(_1862_),
    .Y(_1863_));
 sky130_fd_sc_hd__o32a_1 _4725_ (.A1(_1616_),
    .A2(_0591_),
    .A3(_1855_),
    .B1(_1617_),
    .B2(_0603_),
    .X(_1864_));
 sky130_fd_sc_hd__a21oi_4 _4726_ (.A1(_1610_),
    .A2(_0595_),
    .B1(_1860_),
    .Y(_1865_));
 sky130_fd_sc_hd__a21oi_4 _4727_ (.A1(_1612_),
    .A2(_0598_),
    .B1(_1861_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _4728_ (.A(_1865_),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__nor2_1 _4729_ (.A(\acc3[3] ),
    .B(\acc2[3] ),
    .Y(_1868_));
 sky130_fd_sc_hd__a21oi_2 _4730_ (.A1(\acc3[3] ),
    .A2(\acc2[3] ),
    .B1(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__inv_2 _4731_ (.A(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__o22a_1 _4732_ (.A1(_1626_),
    .A2(_0612_),
    .B1(\acc3[2] ),
    .B2(\acc2[2] ),
    .X(_1871_));
 sky130_fd_sc_hd__inv_2 _4733_ (.A(_1871_),
    .Y(_1872_));
 sky130_fd_sc_hd__a22o_1 _4734_ (.A1(\acc3[1] ),
    .A2(\acc2[1] ),
    .B1(_1628_),
    .B2(_0618_),
    .X(_1873_));
 sky130_fd_sc_hd__or3_1 _4735_ (.A(_1778_),
    .B(_0620_),
    .C(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__o21ai_2 _4736_ (.A1(_1628_),
    .A2(_0618_),
    .B1(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__inv_2 _4737_ (.A(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__o32a_1 _4738_ (.A1(_1635_),
    .A2(_0613_),
    .A3(_1868_),
    .B1(_1636_),
    .B2(_0627_),
    .X(_1877_));
 sky130_fd_sc_hd__o31a_1 _4739_ (.A1(_1870_),
    .A2(_1872_),
    .A3(_1876_),
    .B1(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__or4_4 _4740_ (.A(_1857_),
    .B(_1859_),
    .C(_1867_),
    .D(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__o311a_2 _4741_ (.A1(_1857_),
    .A2(_1859_),
    .A3(_1863_),
    .B1(_1864_),
    .C1(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__a22o_1 _4742_ (.A1(_1579_),
    .A2(_0557_),
    .B1(\acc3[12] ),
    .B2(\acc2[12] ),
    .X(_1881_));
 sky130_fd_sc_hd__o21ai_1 _4743_ (.A1(_1579_),
    .A2(_0557_),
    .B1(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__a22o_1 _4744_ (.A1(_1594_),
    .A2(_0577_),
    .B1(\acc3[8] ),
    .B2(\acc2[8] ),
    .X(_1883_));
 sky130_fd_sc_hd__o21ai_1 _4745_ (.A1(_1594_),
    .A2(_0577_),
    .B1(_1883_),
    .Y(_1884_));
 sky130_fd_sc_hd__a211o_1 _4746_ (.A1(_1643_),
    .A2(_0568_),
    .B1(_1646_),
    .C1(_0572_),
    .X(_1885_));
 sky130_fd_sc_hd__o221a_1 _4747_ (.A1(_1643_),
    .A2(_0568_),
    .B1(_1848_),
    .B2(_1884_),
    .C1(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__o32a_1 _4748_ (.A1(_1649_),
    .A2(_0552_),
    .A3(_1836_),
    .B1(_1650_),
    .B2(_0639_),
    .X(_1887_));
 sky130_fd_sc_hd__o221a_1 _4749_ (.A1(_1839_),
    .A2(_1882_),
    .B1(_1845_),
    .B2(_1886_),
    .C1(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__o31a_2 _4750_ (.A1(_1845_),
    .A2(_1854_),
    .A3(_1880_),
    .B1(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__o22a_1 _4751_ (.A1(_1558_),
    .A2(_0538_),
    .B1(_1654_),
    .B2(_0644_),
    .X(_1890_));
 sky130_fd_sc_hd__inv_2 _4752_ (.A(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__o22a_1 _4753_ (.A1(_1657_),
    .A2(_0648_),
    .B1(\acc3[16] ),
    .B2(\acc2[16] ),
    .X(_1892_));
 sky130_fd_sc_hd__inv_2 _4754_ (.A(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__mux2_2 _4755_ (.A0(_0034_),
    .A1(_0032_),
    .S(_0033_),
    .X(_2370_));
 sky130_fd_sc_hd__mux2_1 _4756_ (.A0(_0001_),
    .A1(_0035_),
    .S(_0033_),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_1 _4757_ (.A0(_0003_),
    .A1(_0002_),
    .S(_0033_),
    .X(_2378_));
 sky130_fd_sc_hd__mux2_1 _4758_ (.A0(_0005_),
    .A1(_0004_),
    .S(_0033_),
    .X(_2379_));
 sky130_fd_sc_hd__mux2_2 _4759_ (.A0(_0007_),
    .A1(_0006_),
    .S(_0033_),
    .X(_2380_));
 sky130_fd_sc_hd__mux2_2 _4760_ (.A0(_0009_),
    .A1(_0008_),
    .S(_0033_),
    .X(_2381_));
 sky130_fd_sc_hd__mux2_2 _4761_ (.A0(_0011_),
    .A1(_0010_),
    .S(_0033_),
    .X(_2382_));
 sky130_fd_sc_hd__mux2_2 _4762_ (.A0(_0013_),
    .A1(_0012_),
    .S(_0033_),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_2 _4763_ (.A0(_0015_),
    .A1(_0014_),
    .S(_0033_),
    .X(_2384_));
 sky130_fd_sc_hd__mux2_1 _4764_ (.A0(_0017_),
    .A1(_0016_),
    .S(_0033_),
    .X(_2385_));
 sky130_fd_sc_hd__mux2_1 _4765_ (.A0(_0019_),
    .A1(_0018_),
    .S(_0033_),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(_0021_),
    .A1(_0020_),
    .S(_0033_),
    .X(_2372_));
 sky130_fd_sc_hd__mux2_2 _4767_ (.A0(_0023_),
    .A1(_0022_),
    .S(_0033_),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_2 _4768_ (.A0(_0025_),
    .A1(_0024_),
    .S(_0033_),
    .X(_2374_));
 sky130_fd_sc_hd__mux2_2 _4769_ (.A0(_0027_),
    .A1(_0026_),
    .S(_0033_),
    .X(_2375_));
 sky130_fd_sc_hd__mux2_1 _4770_ (.A0(_0029_),
    .A1(_0028_),
    .S(_0033_),
    .X(_2376_));
 sky130_fd_sc_hd__mux2_1 _4771_ (.A0(_0030_),
    .A1(_0031_),
    .S(enable),
    .X(_0000_));
 sky130_fd_sc_hd__dfxtp_1 _4772_ (.D(_2370_),
    .Q(net19),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4773_ (.D(_2377_),
    .Q(net26),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4774_ (.D(_2378_),
    .Q(net27),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4775_ (.D(_2379_),
    .Q(net28),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4776_ (.D(_2380_),
    .Q(net29),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4777_ (.D(_2381_),
    .Q(net30),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4778_ (.D(_2382_),
    .Q(net31),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4779_ (.D(_2383_),
    .Q(net32),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4780_ (.D(_2384_),
    .Q(net33),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4781_ (.D(_2385_),
    .Q(net34),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4782_ (.D(_2371_),
    .Q(net20),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4783_ (.D(_2372_),
    .Q(net21),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4784_ (.D(_2373_),
    .Q(net22),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4785_ (.D(_2374_),
    .Q(net23),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4786_ (.D(_2375_),
    .Q(net24),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4787_ (.D(_2376_),
    .Q(net25),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4788_ (.D(_0147_),
    .Q(\acc3[0] ),
    .CLK(_0036_));
 sky130_fd_sc_hd__dfxtp_1 _4789_ (.D(_0148_),
    .Q(\acc3[1] ),
    .CLK(_0037_));
 sky130_fd_sc_hd__dfxtp_1 _4790_ (.D(_0149_),
    .Q(\acc3[2] ),
    .CLK(_0038_));
 sky130_fd_sc_hd__dfxtp_2 _4791_ (.D(_0150_),
    .Q(\acc3[3] ),
    .CLK(_0039_));
 sky130_fd_sc_hd__dfxtp_1 _4792_ (.D(_0151_),
    .Q(\acc3[4] ),
    .CLK(_0040_));
 sky130_fd_sc_hd__dfxtp_1 _4793_ (.D(_0152_),
    .Q(\acc3[5] ),
    .CLK(_0041_));
 sky130_fd_sc_hd__dfxtp_1 _4794_ (.D(_0153_),
    .Q(\acc3[6] ),
    .CLK(_0042_));
 sky130_fd_sc_hd__dfxtp_2 _4795_ (.D(_0154_),
    .Q(\acc3[7] ),
    .CLK(_0043_));
 sky130_fd_sc_hd__dfxtp_1 _4796_ (.D(_0155_),
    .Q(\acc3[8] ),
    .CLK(_0044_));
 sky130_fd_sc_hd__dfxtp_1 _4797_ (.D(_0156_),
    .Q(\acc3[9] ),
    .CLK(_0045_));
 sky130_fd_sc_hd__dfxtp_1 _4798_ (.D(_0157_),
    .Q(\acc3[10] ),
    .CLK(_0046_));
 sky130_fd_sc_hd__dfxtp_1 _4799_ (.D(_0158_),
    .Q(\acc3[11] ),
    .CLK(_0047_));
 sky130_fd_sc_hd__dfxtp_1 _4800_ (.D(_0159_),
    .Q(\acc3[12] ),
    .CLK(_0048_));
 sky130_fd_sc_hd__dfxtp_1 _4801_ (.D(_0160_),
    .Q(\acc3[13] ),
    .CLK(_0049_));
 sky130_fd_sc_hd__dfxtp_1 _4802_ (.D(_0161_),
    .Q(\acc3[14] ),
    .CLK(_0050_));
 sky130_fd_sc_hd__dfxtp_2 _4803_ (.D(_0162_),
    .Q(\acc3[15] ),
    .CLK(_0051_));
 sky130_fd_sc_hd__dfxtp_1 _4804_ (.D(_0163_),
    .Q(\acc3[16] ),
    .CLK(_0052_));
 sky130_fd_sc_hd__dfxtp_1 _4805_ (.D(_0164_),
    .Q(\acc3[17] ),
    .CLK(_0053_));
 sky130_fd_sc_hd__dfxtp_1 _4806_ (.D(_0165_),
    .Q(\acc3[18] ),
    .CLK(_0054_));
 sky130_fd_sc_hd__dfxtp_1 _4807_ (.D(_0166_),
    .Q(\acc3[19] ),
    .CLK(_0055_));
 sky130_fd_sc_hd__dfxtp_1 _4808_ (.D(_0167_),
    .Q(\acc3[20] ),
    .CLK(_0056_));
 sky130_fd_sc_hd__dfxtp_1 _4809_ (.D(_0168_),
    .Q(\acc3[21] ),
    .CLK(_0057_));
 sky130_fd_sc_hd__dfxtp_1 _4810_ (.D(_0169_),
    .Q(\acc3[22] ),
    .CLK(_0058_));
 sky130_fd_sc_hd__dfxtp_2 _4811_ (.D(_0170_),
    .Q(\acc3[23] ),
    .CLK(_0059_));
 sky130_fd_sc_hd__dfxtp_1 _4812_ (.D(_0171_),
    .Q(\acc3[24] ),
    .CLK(_0060_));
 sky130_fd_sc_hd__dfxtp_1 _4813_ (.D(_0172_),
    .Q(\acc3[25] ),
    .CLK(_0061_));
 sky130_fd_sc_hd__dfxtp_1 _4814_ (.D(_0173_),
    .Q(\acc3[26] ),
    .CLK(_0062_));
 sky130_fd_sc_hd__dfxtp_1 _4815_ (.D(_0174_),
    .Q(\acc3[27] ),
    .CLK(_0063_));
 sky130_fd_sc_hd__dfxtp_1 _4816_ (.D(_0175_),
    .Q(\acc3[28] ),
    .CLK(_0064_));
 sky130_fd_sc_hd__dfxtp_1 _4817_ (.D(_0176_),
    .Q(\acc3[29] ),
    .CLK(_0065_));
 sky130_fd_sc_hd__dfxtp_1 _4818_ (.D(_0177_),
    .Q(\acc3[30] ),
    .CLK(_0066_));
 sky130_fd_sc_hd__dfxtp_2 _4819_ (.D(_0178_),
    .Q(\acc3[31] ),
    .CLK(_0067_));
 sky130_fd_sc_hd__dfxtp_1 _4820_ (.D(_0179_),
    .Q(\acc3[32] ),
    .CLK(_0068_));
 sky130_fd_sc_hd__dfxtp_2 _4821_ (.D(_0180_),
    .Q(\acc3[33] ),
    .CLK(_0069_));
 sky130_fd_sc_hd__dfxtp_1 _4822_ (.D(_0181_),
    .Q(\acc3[34] ),
    .CLK(_0070_));
 sky130_fd_sc_hd__dfxtp_2 _4823_ (.D(_0182_),
    .Q(\acc3[35] ),
    .CLK(_0071_));
 sky130_fd_sc_hd__dfxtp_1 _4824_ (.D(_0183_),
    .Q(\acc3[36] ),
    .CLK(_0072_));
 sky130_fd_sc_hd__dfxtp_1 _4825_ (.D(_0184_),
    .Q(net35),
    .CLK(clknet_1_0_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _4826_ (.D(_0185_),
    .Q(\acc3_d2[0] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4827_ (.D(_0186_),
    .Q(\acc3_d2[1] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4828_ (.D(_0187_),
    .Q(\acc3_d2[2] ),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4829_ (.D(_0188_),
    .Q(\acc3_d2[3] ),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_2 _4830_ (.D(_0189_),
    .Q(\acc3_d2[4] ),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4831_ (.D(_0190_),
    .Q(\acc3_d2[5] ),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4832_ (.D(_0191_),
    .Q(\acc3_d2[6] ),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4833_ (.D(_0192_),
    .Q(\acc3_d2[7] ),
    .CLK(word_clk));
 sky130_fd_sc_hd__dfxtp_1 _4834_ (.D(_0193_),
    .Q(\acc3_d2[8] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4835_ (.D(_0194_),
    .Q(\acc3_d2[9] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4836_ (.D(_0195_),
    .Q(\acc3_d2[10] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4837_ (.D(_0196_),
    .Q(\acc3_d2[11] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4838_ (.D(_0197_),
    .Q(\acc3_d2[12] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4839_ (.D(_0198_),
    .Q(\acc3_d2[13] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4840_ (.D(_0199_),
    .Q(\acc3_d2[14] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4841_ (.D(_0200_),
    .Q(\acc3_d2[15] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4842_ (.D(_0201_),
    .Q(\acc3_d2[16] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4843_ (.D(_0202_),
    .Q(\acc3_d2[17] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4844_ (.D(_0203_),
    .Q(\acc3_d2[18] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4845_ (.D(_0204_),
    .Q(\acc3_d2[19] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4846_ (.D(_0205_),
    .Q(\acc3_d2[20] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4847_ (.D(_0206_),
    .Q(\acc3_d2[21] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4848_ (.D(_0207_),
    .Q(\acc3_d2[22] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4849_ (.D(_0208_),
    .Q(\acc3_d2[23] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4850_ (.D(_0209_),
    .Q(\acc3_d2[24] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4851_ (.D(_0210_),
    .Q(\acc3_d2[25] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4852_ (.D(_0211_),
    .Q(\acc3_d2[26] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4853_ (.D(_0212_),
    .Q(\acc3_d2[27] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4854_ (.D(_0213_),
    .Q(\acc3_d2[28] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4855_ (.D(_0214_),
    .Q(\acc3_d2[29] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4856_ (.D(_0215_),
    .Q(\acc3_d2[30] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4857_ (.D(_0216_),
    .Q(\acc3_d2[31] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4858_ (.D(_0217_),
    .Q(\acc3_d2[32] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4859_ (.D(_0218_),
    .Q(\acc3_d2[33] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4860_ (.D(_0219_),
    .Q(\acc3_d2[34] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4861_ (.D(_0220_),
    .Q(\acc3_d2[35] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4862_ (.D(_0221_),
    .Q(\acc3_d2[36] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4863_ (.D(_0222_),
    .Q(\diff1[0] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4864_ (.D(_0223_),
    .Q(\diff1[1] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4865_ (.D(_0224_),
    .Q(\diff1[2] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4866_ (.D(_0225_),
    .Q(\diff1[3] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4867_ (.D(_0226_),
    .Q(\diff1[4] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4868_ (.D(_0227_),
    .Q(\diff1[5] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4869_ (.D(_0228_),
    .Q(\diff1[6] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4870_ (.D(_0229_),
    .Q(\diff1[7] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4871_ (.D(_0230_),
    .Q(\diff1[8] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4872_ (.D(_0231_),
    .Q(\diff1[9] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4873_ (.D(_0232_),
    .Q(\diff1[10] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4874_ (.D(_0233_),
    .Q(\diff1[11] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4875_ (.D(_0234_),
    .Q(\diff1[12] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4876_ (.D(_0235_),
    .Q(\diff1[13] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4877_ (.D(_0236_),
    .Q(\diff1[14] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4878_ (.D(_0237_),
    .Q(\diff1[15] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4879_ (.D(_0238_),
    .Q(\diff1[16] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4880_ (.D(_0239_),
    .Q(\diff1[17] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4881_ (.D(_0240_),
    .Q(\diff1[18] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4882_ (.D(_0241_),
    .Q(\diff1[19] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4883_ (.D(_0242_),
    .Q(\diff1[20] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4884_ (.D(_0243_),
    .Q(\diff1[21] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4885_ (.D(_0244_),
    .Q(\diff1[22] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4886_ (.D(_0245_),
    .Q(\diff1[23] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4887_ (.D(_0246_),
    .Q(\diff1[24] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4888_ (.D(_0247_),
    .Q(\diff1[25] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4889_ (.D(_0248_),
    .Q(\diff1[26] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4890_ (.D(_0249_),
    .Q(\diff1[27] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4891_ (.D(_0250_),
    .Q(\diff1[28] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4892_ (.D(_0251_),
    .Q(\diff1[29] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4893_ (.D(_0252_),
    .Q(\diff1[30] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4894_ (.D(_0253_),
    .Q(\diff1[31] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4895_ (.D(_0254_),
    .Q(\diff1[32] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4896_ (.D(_0255_),
    .Q(\diff1[33] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4897_ (.D(_0256_),
    .Q(\diff1[34] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4898_ (.D(_0257_),
    .Q(\diff1[35] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4899_ (.D(_0258_),
    .Q(\diff1[36] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4900_ (.D(_0259_),
    .Q(\diff2[0] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4901_ (.D(_0260_),
    .Q(\diff2[1] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4902_ (.D(_0261_),
    .Q(\diff2[2] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4903_ (.D(_0262_),
    .Q(\diff2[3] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4904_ (.D(_0263_),
    .Q(\diff2[4] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4905_ (.D(_0264_),
    .Q(\diff2[5] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4906_ (.D(_0265_),
    .Q(\diff2[6] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4907_ (.D(_0266_),
    .Q(\diff2[7] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4908_ (.D(_0267_),
    .Q(\diff2[8] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4909_ (.D(_0268_),
    .Q(\diff2[9] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4910_ (.D(_0269_),
    .Q(\diff2[10] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4911_ (.D(_0270_),
    .Q(\diff2[11] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4912_ (.D(_0271_),
    .Q(\diff2[12] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4913_ (.D(_0272_),
    .Q(\diff2[13] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4914_ (.D(_0273_),
    .Q(\diff2[14] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4915_ (.D(_0274_),
    .Q(\diff2[15] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4916_ (.D(_0275_),
    .Q(\diff2[16] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4917_ (.D(_0276_),
    .Q(\diff2[17] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4918_ (.D(_0277_),
    .Q(\diff2[18] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4919_ (.D(_0278_),
    .Q(\diff2[19] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4920_ (.D(_0279_),
    .Q(\diff2[20] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4921_ (.D(_0280_),
    .Q(\diff2[21] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4922_ (.D(_0281_),
    .Q(\diff2[22] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4923_ (.D(_0282_),
    .Q(\diff2[23] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4924_ (.D(_0283_),
    .Q(\diff2[24] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4925_ (.D(_0284_),
    .Q(\diff2[25] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4926_ (.D(_0285_),
    .Q(\diff2[26] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4927_ (.D(_0286_),
    .Q(\diff2[27] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4928_ (.D(_0287_),
    .Q(\diff2[28] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4929_ (.D(_0288_),
    .Q(\diff2[29] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4930_ (.D(_0289_),
    .Q(\diff2[30] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4931_ (.D(_0290_),
    .Q(\diff2[31] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4932_ (.D(_0291_),
    .Q(\diff2[32] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4933_ (.D(_0292_),
    .Q(\diff2[33] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4934_ (.D(_0293_),
    .Q(\diff2[34] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4935_ (.D(_0294_),
    .Q(\diff2[35] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4936_ (.D(_0295_),
    .Q(\diff2[36] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4937_ (.D(_0296_),
    .Q(\diff3[0] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4938_ (.D(_0297_),
    .Q(\diff3[1] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4939_ (.D(_0298_),
    .Q(\diff3[2] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4940_ (.D(_0299_),
    .Q(\diff3[3] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4941_ (.D(_0300_),
    .Q(\diff3[4] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_2 _4942_ (.D(_0301_),
    .Q(\diff3[5] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4943_ (.D(_0302_),
    .Q(\diff3[6] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4944_ (.D(_0303_),
    .Q(\diff3[7] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4945_ (.D(_0304_),
    .Q(\diff3[8] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4946_ (.D(_0305_),
    .Q(\diff3[9] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4947_ (.D(_0306_),
    .Q(\diff3[10] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4948_ (.D(_0307_),
    .Q(\diff3[11] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4949_ (.D(_0308_),
    .Q(\diff3[12] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4950_ (.D(_0309_),
    .Q(\diff3[13] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4951_ (.D(_0310_),
    .Q(\diff3[14] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4952_ (.D(_0311_),
    .Q(\diff3[15] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4953_ (.D(_0312_),
    .Q(\diff3[16] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4954_ (.D(_0313_),
    .Q(\diff3[17] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4955_ (.D(_0314_),
    .Q(\diff3[18] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4956_ (.D(_0315_),
    .Q(\diff3[19] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4957_ (.D(_0316_),
    .Q(\diff3[20] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4958_ (.D(_0317_),
    .Q(\diff3[21] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4959_ (.D(_0318_),
    .Q(\diff3[22] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4960_ (.D(_0319_),
    .Q(\diff3[23] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4961_ (.D(_0320_),
    .Q(\diff3[24] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4962_ (.D(_0321_),
    .Q(\diff3[25] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4963_ (.D(_0322_),
    .Q(\diff3[26] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4964_ (.D(_0323_),
    .Q(\diff3[27] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4965_ (.D(_0324_),
    .Q(\diff3[28] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4966_ (.D(_0325_),
    .Q(\diff3[29] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4967_ (.D(_0326_),
    .Q(\diff3[30] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4968_ (.D(_0327_),
    .Q(\diff3[31] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4969_ (.D(_0328_),
    .Q(\diff3[32] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4970_ (.D(_0329_),
    .Q(\diff3[33] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4971_ (.D(_0330_),
    .Q(\diff3[34] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4972_ (.D(_0331_),
    .Q(\diff3[35] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4973_ (.D(_0332_),
    .Q(\diff3[36] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4974_ (.D(_0333_),
    .Q(\diff1_d[0] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4975_ (.D(_0334_),
    .Q(\diff1_d[1] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4976_ (.D(_0335_),
    .Q(\diff1_d[2] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4977_ (.D(_0336_),
    .Q(\diff1_d[3] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_2 _4978_ (.D(_0337_),
    .Q(\diff1_d[4] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4979_ (.D(_0338_),
    .Q(\diff1_d[5] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4980_ (.D(_0339_),
    .Q(\diff1_d[6] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4981_ (.D(_0340_),
    .Q(\diff1_d[7] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _4982_ (.D(_0341_),
    .Q(\diff1_d[8] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4983_ (.D(_0342_),
    .Q(\diff1_d[9] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4984_ (.D(_0343_),
    .Q(\diff1_d[10] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4985_ (.D(_0344_),
    .Q(\diff1_d[11] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4986_ (.D(_0345_),
    .Q(\diff1_d[12] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4987_ (.D(_0346_),
    .Q(\diff1_d[13] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4988_ (.D(_0347_),
    .Q(\diff1_d[14] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4989_ (.D(_0348_),
    .Q(\diff1_d[15] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4990_ (.D(_0349_),
    .Q(\diff1_d[16] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4991_ (.D(_0350_),
    .Q(\diff1_d[17] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4992_ (.D(_0351_),
    .Q(\diff1_d[18] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4993_ (.D(_0352_),
    .Q(\diff1_d[19] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4994_ (.D(_0353_),
    .Q(\diff1_d[20] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4995_ (.D(_0354_),
    .Q(\diff1_d[21] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4996_ (.D(_0355_),
    .Q(\diff1_d[22] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4997_ (.D(_0356_),
    .Q(\diff1_d[23] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _4998_ (.D(_0357_),
    .Q(\diff1_d[24] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _4999_ (.D(_0358_),
    .Q(\diff1_d[25] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5000_ (.D(_0359_),
    .Q(\diff1_d[26] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5001_ (.D(_0360_),
    .Q(\diff1_d[27] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5002_ (.D(_0361_),
    .Q(\diff1_d[28] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5003_ (.D(_0362_),
    .Q(\diff1_d[29] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5004_ (.D(_0363_),
    .Q(\diff1_d[30] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5005_ (.D(_0364_),
    .Q(\diff1_d[31] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5006_ (.D(_0365_),
    .Q(\diff1_d[32] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5007_ (.D(_0366_),
    .Q(\diff1_d[33] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5008_ (.D(_0367_),
    .Q(\diff1_d[34] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5009_ (.D(_0368_),
    .Q(\diff1_d[35] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5010_ (.D(_0369_),
    .Q(\diff1_d[36] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5011_ (.D(_0370_),
    .Q(\diff2_d[0] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _5012_ (.D(_0371_),
    .Q(\diff2_d[1] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _5013_ (.D(_0372_),
    .Q(\diff2_d[2] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _5014_ (.D(_0373_),
    .Q(\diff2_d[3] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_2 _5015_ (.D(_0374_),
    .Q(\diff2_d[4] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _5016_ (.D(_0375_),
    .Q(\diff2_d[5] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _5017_ (.D(_0376_),
    .Q(\diff2_d[6] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _5018_ (.D(_0377_),
    .Q(\diff2_d[7] ),
    .CLK(net38));
 sky130_fd_sc_hd__dfxtp_1 _5019_ (.D(_0378_),
    .Q(\diff2_d[8] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5020_ (.D(_0379_),
    .Q(\diff2_d[9] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5021_ (.D(_0380_),
    .Q(\diff2_d[10] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5022_ (.D(_0381_),
    .Q(\diff2_d[11] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5023_ (.D(_0382_),
    .Q(\diff2_d[12] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5024_ (.D(_0383_),
    .Q(\diff2_d[13] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5025_ (.D(_0384_),
    .Q(\diff2_d[14] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5026_ (.D(_0385_),
    .Q(\diff2_d[15] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5027_ (.D(_0386_),
    .Q(\diff2_d[16] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5028_ (.D(_0387_),
    .Q(\diff2_d[17] ),
    .CLK(net37));
 sky130_fd_sc_hd__dfxtp_1 _5029_ (.D(_0388_),
    .Q(\diff2_d[18] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5030_ (.D(_0389_),
    .Q(\diff2_d[19] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5031_ (.D(_0390_),
    .Q(\diff2_d[20] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5032_ (.D(_0391_),
    .Q(\diff2_d[21] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5033_ (.D(_0392_),
    .Q(\diff2_d[22] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5034_ (.D(_0393_),
    .Q(\diff2_d[23] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5035_ (.D(_0394_),
    .Q(\diff2_d[24] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5036_ (.D(_0395_),
    .Q(\diff2_d[25] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5037_ (.D(_0396_),
    .Q(\diff2_d[26] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5038_ (.D(_0397_),
    .Q(\diff2_d[27] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5039_ (.D(_0398_),
    .Q(\diff2_d[28] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5040_ (.D(_0399_),
    .Q(\diff2_d[29] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5041_ (.D(_0400_),
    .Q(\diff2_d[30] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5042_ (.D(_0401_),
    .Q(\diff2_d[31] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5043_ (.D(_0402_),
    .Q(\diff2_d[32] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5044_ (.D(_0403_),
    .Q(\diff2_d[33] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5045_ (.D(_0404_),
    .Q(\diff2_d[34] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5046_ (.D(_0405_),
    .Q(\diff2_d[35] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5047_ (.D(_0406_),
    .Q(\diff2_d[36] ),
    .CLK(net36));
 sky130_fd_sc_hd__dfxtp_1 _5048_ (.D(_0407_),
    .Q(\word_count[0] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5049_ (.D(_0408_),
    .Q(\word_count[1] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5050_ (.D(_0409_),
    .Q(\word_count[2] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5051_ (.D(_0410_),
    .Q(\word_count[3] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5052_ (.D(_0411_),
    .Q(\word_count[4] ),
    .CLK(clknet_1_0_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5053_ (.D(_0412_),
    .Q(\word_count[5] ),
    .CLK(clknet_1_0_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5054_ (.D(_0413_),
    .Q(\word_count[6] ),
    .CLK(clknet_1_0_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5055_ (.D(_0414_),
    .Q(\word_count[7] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5056_ (.D(_0415_),
    .Q(\word_count[8] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5057_ (.D(_0416_),
    .Q(\word_count[9] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5058_ (.D(_0417_),
    .Q(\word_count[10] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5059_ (.D(_0418_),
    .Q(\word_count[11] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_2 _5060_ (.D(_0419_),
    .Q(\word_count[12] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5061_ (.D(_0420_),
    .Q(\word_count[13] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5062_ (.D(_0421_),
    .Q(\word_count[14] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5063_ (.D(_0422_),
    .Q(\word_count[15] ),
    .CLK(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dfxtp_1 _5064_ (.D(_0423_),
    .Q(\acc1[0] ),
    .CLK(_0073_));
 sky130_fd_sc_hd__dfxtp_1 _5065_ (.D(_0424_),
    .Q(\acc1[1] ),
    .CLK(_0074_));
 sky130_fd_sc_hd__dfxtp_1 _5066_ (.D(_0425_),
    .Q(\acc1[2] ),
    .CLK(_0075_));
 sky130_fd_sc_hd__dfxtp_1 _5067_ (.D(_0426_),
    .Q(\acc1[3] ),
    .CLK(_0076_));
 sky130_fd_sc_hd__dfxtp_1 _5068_ (.D(_0427_),
    .Q(\acc1[4] ),
    .CLK(_0077_));
 sky130_fd_sc_hd__dfxtp_1 _5069_ (.D(_0428_),
    .Q(\acc1[5] ),
    .CLK(_0078_));
 sky130_fd_sc_hd__dfxtp_1 _5070_ (.D(_0429_),
    .Q(\acc1[6] ),
    .CLK(_0079_));
 sky130_fd_sc_hd__dfxtp_1 _5071_ (.D(_0430_),
    .Q(\acc1[7] ),
    .CLK(_0080_));
 sky130_fd_sc_hd__dfxtp_1 _5072_ (.D(_0431_),
    .Q(\acc1[8] ),
    .CLK(_0081_));
 sky130_fd_sc_hd__dfxtp_1 _5073_ (.D(_0432_),
    .Q(\acc1[9] ),
    .CLK(_0082_));
 sky130_fd_sc_hd__dfxtp_1 _5074_ (.D(_0433_),
    .Q(\acc1[10] ),
    .CLK(_0083_));
 sky130_fd_sc_hd__dfxtp_1 _5075_ (.D(_0434_),
    .Q(\acc1[11] ),
    .CLK(_0084_));
 sky130_fd_sc_hd__dfxtp_1 _5076_ (.D(_0435_),
    .Q(\acc1[12] ),
    .CLK(_0085_));
 sky130_fd_sc_hd__dfxtp_1 _5077_ (.D(_0436_),
    .Q(\acc1[13] ),
    .CLK(_0086_));
 sky130_fd_sc_hd__dfxtp_1 _5078_ (.D(_0437_),
    .Q(\acc1[14] ),
    .CLK(_0087_));
 sky130_fd_sc_hd__dfxtp_1 _5079_ (.D(_0438_),
    .Q(\acc1[15] ),
    .CLK(_0088_));
 sky130_fd_sc_hd__dfxtp_1 _5080_ (.D(_0439_),
    .Q(\acc1[16] ),
    .CLK(_0089_));
 sky130_fd_sc_hd__dfxtp_1 _5081_ (.D(_0440_),
    .Q(\acc1[17] ),
    .CLK(_0090_));
 sky130_fd_sc_hd__dfxtp_1 _5082_ (.D(_0441_),
    .Q(\acc1[18] ),
    .CLK(_0091_));
 sky130_fd_sc_hd__dfxtp_1 _5083_ (.D(_0442_),
    .Q(\acc1[19] ),
    .CLK(_0092_));
 sky130_fd_sc_hd__dfxtp_1 _5084_ (.D(_0443_),
    .Q(\acc1[20] ),
    .CLK(_0093_));
 sky130_fd_sc_hd__dfxtp_1 _5085_ (.D(_0444_),
    .Q(\acc1[21] ),
    .CLK(_0094_));
 sky130_fd_sc_hd__dfxtp_1 _5086_ (.D(_0445_),
    .Q(\acc1[22] ),
    .CLK(_0095_));
 sky130_fd_sc_hd__dfxtp_1 _5087_ (.D(_0446_),
    .Q(\acc1[23] ),
    .CLK(_0096_));
 sky130_fd_sc_hd__dfxtp_1 _5088_ (.D(_0447_),
    .Q(\acc1[24] ),
    .CLK(_0097_));
 sky130_fd_sc_hd__dfxtp_1 _5089_ (.D(_0448_),
    .Q(\acc1[25] ),
    .CLK(_0098_));
 sky130_fd_sc_hd__dfxtp_2 _5090_ (.D(_0449_),
    .Q(\acc1[26] ),
    .CLK(_0099_));
 sky130_fd_sc_hd__dfxtp_1 _5091_ (.D(_0450_),
    .Q(\acc1[27] ),
    .CLK(_0100_));
 sky130_fd_sc_hd__dfxtp_1 _5092_ (.D(_0451_),
    .Q(\acc1[28] ),
    .CLK(_0101_));
 sky130_fd_sc_hd__dfxtp_1 _5093_ (.D(_0452_),
    .Q(\acc1[29] ),
    .CLK(_0102_));
 sky130_fd_sc_hd__dfxtp_1 _5094_ (.D(_0453_),
    .Q(\acc1[30] ),
    .CLK(_0103_));
 sky130_fd_sc_hd__dfxtp_1 _5095_ (.D(_0454_),
    .Q(\acc1[31] ),
    .CLK(_0104_));
 sky130_fd_sc_hd__dfxtp_1 _5096_ (.D(_0455_),
    .Q(\acc1[32] ),
    .CLK(_0105_));
 sky130_fd_sc_hd__dfxtp_1 _5097_ (.D(_0456_),
    .Q(\acc1[33] ),
    .CLK(_0106_));
 sky130_fd_sc_hd__dfxtp_1 _5098_ (.D(_0457_),
    .Q(\acc1[34] ),
    .CLK(_0107_));
 sky130_fd_sc_hd__dfxtp_1 _5099_ (.D(_0458_),
    .Q(\acc1[35] ),
    .CLK(_0108_));
 sky130_fd_sc_hd__dfxtp_1 _5100_ (.D(_0459_),
    .Q(\acc1[36] ),
    .CLK(_0109_));
 sky130_fd_sc_hd__dfxtp_1 _5101_ (.D(_0460_),
    .Q(\acc2[0] ),
    .CLK(_0110_));
 sky130_fd_sc_hd__dfxtp_1 _5102_ (.D(_0461_),
    .Q(\acc2[1] ),
    .CLK(_0111_));
 sky130_fd_sc_hd__dfxtp_1 _5103_ (.D(_0462_),
    .Q(\acc2[2] ),
    .CLK(_0112_));
 sky130_fd_sc_hd__dfxtp_2 _5104_ (.D(_0463_),
    .Q(\acc2[3] ),
    .CLK(_0113_));
 sky130_fd_sc_hd__dfxtp_1 _5105_ (.D(_0464_),
    .Q(\acc2[4] ),
    .CLK(_0114_));
 sky130_fd_sc_hd__dfxtp_1 _5106_ (.D(_0465_),
    .Q(\acc2[5] ),
    .CLK(_0115_));
 sky130_fd_sc_hd__dfxtp_1 _5107_ (.D(_0466_),
    .Q(\acc2[6] ),
    .CLK(_0116_));
 sky130_fd_sc_hd__dfxtp_2 _5108_ (.D(_0467_),
    .Q(\acc2[7] ),
    .CLK(_0117_));
 sky130_fd_sc_hd__dfxtp_1 _5109_ (.D(_0468_),
    .Q(\acc2[8] ),
    .CLK(_0118_));
 sky130_fd_sc_hd__dfxtp_1 _5110_ (.D(_0469_),
    .Q(\acc2[9] ),
    .CLK(_0119_));
 sky130_fd_sc_hd__dfxtp_1 _5111_ (.D(_0470_),
    .Q(\acc2[10] ),
    .CLK(_0120_));
 sky130_fd_sc_hd__dfxtp_1 _5112_ (.D(_0471_),
    .Q(\acc2[11] ),
    .CLK(_0121_));
 sky130_fd_sc_hd__dfxtp_1 _5113_ (.D(_0472_),
    .Q(\acc2[12] ),
    .CLK(_0122_));
 sky130_fd_sc_hd__dfxtp_1 _5114_ (.D(_0473_),
    .Q(\acc2[13] ),
    .CLK(_0123_));
 sky130_fd_sc_hd__dfxtp_1 _5115_ (.D(_0474_),
    .Q(\acc2[14] ),
    .CLK(_0124_));
 sky130_fd_sc_hd__dfxtp_2 _5116_ (.D(_0475_),
    .Q(\acc2[15] ),
    .CLK(_0125_));
 sky130_fd_sc_hd__dfxtp_1 _5117_ (.D(_0476_),
    .Q(\acc2[16] ),
    .CLK(_0126_));
 sky130_fd_sc_hd__dfxtp_1 _5118_ (.D(_0477_),
    .Q(\acc2[17] ),
    .CLK(_0127_));
 sky130_fd_sc_hd__dfxtp_1 _5119_ (.D(_0478_),
    .Q(\acc2[18] ),
    .CLK(_0128_));
 sky130_fd_sc_hd__dfxtp_1 _5120_ (.D(_0479_),
    .Q(\acc2[19] ),
    .CLK(_0129_));
 sky130_fd_sc_hd__dfxtp_1 _5121_ (.D(_0480_),
    .Q(\acc2[20] ),
    .CLK(_0130_));
 sky130_fd_sc_hd__dfxtp_1 _5122_ (.D(_0481_),
    .Q(\acc2[21] ),
    .CLK(_0131_));
 sky130_fd_sc_hd__dfxtp_1 _5123_ (.D(_0482_),
    .Q(\acc2[22] ),
    .CLK(_0132_));
 sky130_fd_sc_hd__dfxtp_2 _5124_ (.D(_0483_),
    .Q(\acc2[23] ),
    .CLK(_0133_));
 sky130_fd_sc_hd__dfxtp_1 _5125_ (.D(_0484_),
    .Q(\acc2[24] ),
    .CLK(_0134_));
 sky130_fd_sc_hd__dfxtp_1 _5126_ (.D(_0485_),
    .Q(\acc2[25] ),
    .CLK(_0135_));
 sky130_fd_sc_hd__dfxtp_1 _5127_ (.D(_0486_),
    .Q(\acc2[26] ),
    .CLK(_0136_));
 sky130_fd_sc_hd__dfxtp_1 _5128_ (.D(_0487_),
    .Q(\acc2[27] ),
    .CLK(_0137_));
 sky130_fd_sc_hd__dfxtp_1 _5129_ (.D(_0488_),
    .Q(\acc2[28] ),
    .CLK(_0138_));
 sky130_fd_sc_hd__dfxtp_1 _5130_ (.D(_0489_),
    .Q(\acc2[29] ),
    .CLK(_0139_));
 sky130_fd_sc_hd__dfxtp_1 _5131_ (.D(_0490_),
    .Q(\acc2[30] ),
    .CLK(_0140_));
 sky130_fd_sc_hd__dfxtp_2 _5132_ (.D(_0491_),
    .Q(\acc2[31] ),
    .CLK(_0141_));
 sky130_fd_sc_hd__dfxtp_1 _5133_ (.D(_0492_),
    .Q(\acc2[32] ),
    .CLK(_0142_));
 sky130_fd_sc_hd__dfxtp_2 _5134_ (.D(_0493_),
    .Q(\acc2[33] ),
    .CLK(_0143_));
 sky130_fd_sc_hd__dfxtp_1 _5135_ (.D(_0494_),
    .Q(\acc2[34] ),
    .CLK(_0144_));
 sky130_fd_sc_hd__dfxtp_2 _5136_ (.D(_0495_),
    .Q(\acc2[35] ),
    .CLK(_0145_));
 sky130_fd_sc_hd__dfxtp_1 _5137_ (.D(_0496_),
    .Q(\acc2[36] ),
    .CLK(_0146_));
 sky130_fd_sc_hd__dfxtp_1 _5138_ (.D(_0497_),
    .Q(enable),
    .CLK(clknet_1_0_0_mclk1));
 sky130_fd_sc_hd__dfxtp_4 _5139_ (.D(_0498_),
    .Q(word_clk),
    .CLK(clknet_1_0_0_mclk1));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(dec_rate[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dec_rate[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(dec_rate[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(dec_rate[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(dec_rate[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(dec_rate[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(dec_rate[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(dec_rate[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(dec_rate[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(dec_rate[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(dec_rate[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(dec_rate[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(dec_rate[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(dec_rate[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(dec_rate[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(dec_rate[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(mdata1),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(reset),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 output19 (.A(net19),
    .X(DATA[0]));
 sky130_fd_sc_hd__clkbuf_2 output20 (.A(net20),
    .X(DATA[10]));
 sky130_fd_sc_hd__clkbuf_2 output21 (.A(net21),
    .X(DATA[11]));
 sky130_fd_sc_hd__clkbuf_2 output22 (.A(net22),
    .X(DATA[12]));
 sky130_fd_sc_hd__clkbuf_2 output23 (.A(net23),
    .X(DATA[13]));
 sky130_fd_sc_hd__clkbuf_2 output24 (.A(net24),
    .X(DATA[14]));
 sky130_fd_sc_hd__clkbuf_2 output25 (.A(net25),
    .X(DATA[15]));
 sky130_fd_sc_hd__clkbuf_2 output26 (.A(net26),
    .X(DATA[1]));
 sky130_fd_sc_hd__clkbuf_2 output27 (.A(net27),
    .X(DATA[2]));
 sky130_fd_sc_hd__clkbuf_2 output28 (.A(net28),
    .X(DATA[3]));
 sky130_fd_sc_hd__clkbuf_2 output29 (.A(net29),
    .X(DATA[4]));
 sky130_fd_sc_hd__clkbuf_2 output30 (.A(net30),
    .X(DATA[5]));
 sky130_fd_sc_hd__clkbuf_2 output31 (.A(net31),
    .X(DATA[6]));
 sky130_fd_sc_hd__clkbuf_2 output32 (.A(net32),
    .X(DATA[7]));
 sky130_fd_sc_hd__clkbuf_2 output33 (.A(net33),
    .X(DATA[8]));
 sky130_fd_sc_hd__clkbuf_2 output34 (.A(net34),
    .X(DATA[9]));
 sky130_fd_sc_hd__clkbuf_2 output35 (.A(net35),
    .X(data_en));
 sky130_fd_sc_hd__clkbuf_16 repeater36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_16 repeater37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_16 repeater38 (.A(word_clk),
    .X(net38));
 sky130_fd_sc_hd__inv_2 _2926__1 (.A(clknet_1_0_0_mclk1),
    .Y(net39));
 sky130_fd_sc_hd__inv_2 _2926__2 (.A(clknet_1_0_0_mclk1),
    .Y(net40));
 sky130_fd_sc_hd__inv_2 _2926__3 (.A(clknet_1_0_0_mclk1),
    .Y(net41));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_mclk1 (.A(clknet_0_mclk1),
    .X(clknet_1_0_0_mclk1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_mclk1 (.A(clknet_0_mclk1),
    .X(clknet_1_1_0_mclk1));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(net95),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net96),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(_0776_),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_0776_),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_0776_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(_0776_),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(_0803_),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(_0803_),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(_0798_),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(_0779_),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(_0779_),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(_0809_),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(_0809_),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(_0801_),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(_0801_),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer16 (.A(_0793_),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(_0793_),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(_0805_),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(_0805_),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer20 (.A(_0795_),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(_0795_),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer22 (.A(_0797_),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(_0797_),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(_0781_),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer25 (.A(_0781_),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(_0785_),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer27 (.A(_0785_),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(_0807_),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer29 (.A(_0791_),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(_0791_),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer31 (.A(_0783_),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer32 (.A(_0783_),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer33 (.A(_0788_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(_0787_),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(_0787_),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(_0790_),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(_0800_),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(_0799_),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(_0799_),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(_0806_),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(_0780_),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(_0792_),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(_0782_),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net17),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(_0784_),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(_0789_),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(_0789_),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer48 (.A(_0802_),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(_0804_),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(_0796_),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(_0786_),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(_0794_),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(_0808_),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(_0778_),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(_0778_),
    .X(net96));
endmodule
