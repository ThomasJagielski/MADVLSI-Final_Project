magic
tech sky130A
magscale 1 2
timestamp 1619963145
<< obsli1 >>
rect 1104 2159 14168 15249
<< obsm1 >>
rect 474 2128 14168 15280
<< metal2 >>
rect 3698 16635 3754 17435
rect 11058 16635 11114 17435
rect 478 0 534 800
rect 7838 0 7894 800
<< obsm2 >>
rect 480 16579 3642 16635
rect 3810 16579 11002 16635
rect 11170 16579 13506 16635
rect 480 856 13506 16579
rect 590 711 7782 856
rect 7950 711 13506 856
<< metal3 >>
rect 14491 11568 15291 11688
rect 0 10888 800 11008
rect 14491 688 15291 808
<< obsm3 >>
rect 800 11768 14491 15265
rect 800 11488 14411 11768
rect 800 11088 14491 11488
rect 880 10808 14491 11088
rect 800 888 14491 10808
rect 800 715 14411 888
<< metal4 >>
rect 3121 2128 3441 15280
rect 5299 2128 5619 15280
rect 7476 2128 7796 15280
rect 9653 2128 9973 15280
rect 11831 2128 12151 15280
<< obsm4 >>
rect 5699 2128 7396 15280
rect 7876 2128 9573 15280
rect 10053 2128 11751 15280
<< metal5 >>
rect 1104 12848 14168 13168
rect 1104 10672 14168 10992
rect 1104 8496 14168 8816
rect 1104 6320 14168 6640
rect 1104 4144 14168 4464
<< labels >>
rlabel metal2 s 11058 16635 11114 17435 6 clk
port 1 nsew signal input
rlabel metal2 s 478 0 534 800 6 counter[0]
port 2 nsew signal output
rlabel metal3 s 14491 688 15291 808 6 counter[1]
port 3 nsew signal output
rlabel metal3 s 14491 11568 15291 11688 6 counter[2]
port 4 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 counter[3]
port 5 nsew signal output
rlabel metal2 s 3698 16635 3754 17435 6 counter[4]
port 6 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 counter[5]
port 7 nsew signal output
rlabel metal4 s 11831 2128 12151 15280 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 7476 2128 7796 15280 6 VPWR
port 9 nsew power bidirectional
rlabel metal4 s 3121 2128 3441 15280 6 VPWR
port 10 nsew power bidirectional
rlabel metal5 s 1104 12848 14168 13168 6 VPWR
port 11 nsew power bidirectional
rlabel metal5 s 1104 8496 14168 8816 6 VPWR
port 12 nsew power bidirectional
rlabel metal5 s 1104 4144 14168 4464 6 VPWR
port 13 nsew power bidirectional
rlabel metal4 s 9653 2128 9973 15280 6 VGND
port 14 nsew ground bidirectional
rlabel metal4 s 5299 2128 5619 15280 6 VGND
port 15 nsew ground bidirectional
rlabel metal5 s 1104 10672 14168 10992 6 VGND
port 16 nsew ground bidirectional
rlabel metal5 s 1104 6320 14168 6640 6 VGND
port 17 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 15291 17435
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/counter/runs/02-05_13-40/results/magic/counter.gds
string GDS_END 237926
string GDS_START 96820
<< end >>

