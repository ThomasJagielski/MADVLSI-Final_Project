magic
tech sky130A
timestamp 1620753533
<< poly >>
rect -85 3505 -45 3515
rect -85 3485 -75 3505
rect -55 3485 -45 3505
rect -85 3475 -45 3485
rect -85 3040 -65 3475
rect 17815 3345 17855 3355
rect 17815 3325 17825 3345
rect 17845 3325 17855 3345
rect -85 3030 -45 3040
rect -85 3010 -75 3030
rect -55 3010 -45 3030
rect -85 3000 -45 3010
rect 17815 3000 17855 3325
rect 17815 2990 18005 3000
rect 17815 2975 17975 2990
rect 17965 2970 17975 2975
rect 17995 2970 18005 2990
rect 17965 2960 18005 2970
rect 8780 1505 8825 1515
rect 8780 1485 8790 1505
rect 8815 1485 8825 1505
rect 8780 1475 8825 1485
rect 26820 1465 26865 1475
rect 26820 1445 26830 1465
rect 26855 1445 26865 1465
rect 26820 1435 26865 1445
rect 8785 -1760 8830 -1750
rect 8785 -1780 8795 -1760
rect 8820 -1780 8830 -1760
rect 8785 -1790 8830 -1780
rect 26820 -1800 26865 -1790
rect 26820 -1820 26830 -1800
rect 26855 -1820 26865 -1800
rect 26820 -1830 26865 -1820
rect -85 -2000 -35 -1985
rect -85 -2020 -70 -2000
rect -50 -2020 -35 -2000
rect -85 -2125 -35 -2020
rect -85 -2145 -70 -2125
rect -50 -2145 -35 -2125
rect -85 -2160 -35 -2145
rect 17955 -2040 18005 -2025
rect 17955 -2060 17970 -2040
rect 17990 -2060 18005 -2040
rect 17955 -2165 18005 -2060
rect 17955 -2185 17970 -2165
rect 17990 -2185 18005 -2165
rect 17955 -2200 18005 -2185
rect 17615 -2555 17965 -2545
rect 17615 -2560 17930 -2555
rect 17615 -2580 17625 -2560
rect 17645 -2580 17930 -2560
rect 17955 -2580 17965 -2555
rect 17615 -2590 17965 -2580
<< polycont >>
rect -75 3485 -55 3505
rect 17825 3325 17845 3345
rect -75 3010 -55 3030
rect 17975 2970 17995 2990
rect 8790 1485 8815 1505
rect 26830 1445 26855 1465
rect 8795 -1780 8820 -1760
rect 26830 -1820 26855 -1800
rect -70 -2020 -50 -2000
rect -70 -2145 -50 -2125
rect 17970 -2060 17990 -2040
rect 17970 -2185 17990 -2165
rect 17625 -2580 17645 -2560
rect 17930 -2580 17955 -2555
<< locali >>
rect -165 5420 17905 5460
rect -165 3425 -135 5420
rect -85 5320 17855 5360
rect -85 3505 -45 5320
rect -85 3485 -75 3505
rect -55 3485 -45 3505
rect -85 3475 -45 3485
rect -165 3390 55 3425
rect -165 -2055 -135 3390
rect 17815 3345 17855 5320
rect 17815 3325 17825 3345
rect 17845 3325 17855 3345
rect 17815 3315 17855 3325
rect 17875 3385 17905 5420
rect 17875 3350 18095 3385
rect -85 3030 35 3040
rect -85 3010 -75 3030
rect -55 3010 35 3030
rect -85 3000 35 3010
rect -75 -1985 -45 3000
rect 8780 1505 8825 1515
rect 8780 1485 8790 1505
rect 8815 1485 8825 1505
rect 8780 1475 8825 1485
rect 8980 1285 9085 1305
rect 8980 1215 9000 1285
rect 9065 1215 9085 1285
rect 8980 1180 9085 1215
rect 7345 1140 9085 1180
rect 7440 1100 7480 1110
rect 7290 1080 7450 1100
rect 7470 1080 7480 1100
rect 7290 1060 7480 1080
rect 8980 -385 9085 1140
rect 8980 -405 9260 -385
rect 17550 -1310 17610 -1300
rect 17550 -1325 17560 -1310
rect 15870 -1350 17560 -1325
rect 17600 -1350 17610 -1310
rect 17550 -1360 17610 -1350
rect 8600 -1435 9180 -1425
rect 8600 -1455 8610 -1435
rect 8630 -1455 9150 -1435
rect 9170 -1455 9180 -1435
rect 8600 -1465 9180 -1455
rect 8785 -1760 8830 -1750
rect 8785 -1780 8795 -1760
rect 8820 -1780 8830 -1760
rect 8785 -1790 8830 -1780
rect -85 -2000 -35 -1985
rect -85 -2020 -70 -2000
rect -50 -2020 -35 -2000
rect -85 -2035 -35 -2020
rect -165 -2090 65 -2055
rect 17875 -2095 17905 3350
rect 17965 2990 18075 3000
rect 17965 2970 17975 2990
rect 17995 2970 18075 2990
rect 17965 2960 18075 2970
rect 17965 -2025 17995 2960
rect 26820 1465 26865 1475
rect 26820 1445 26830 1465
rect 26855 1445 26865 1465
rect 26820 1435 26865 1445
rect 27020 1245 27125 1265
rect 27020 1175 27040 1245
rect 27105 1175 27125 1245
rect 27020 1140 27125 1175
rect 25385 1100 27125 1140
rect 25330 1050 25520 1060
rect 25330 1030 25490 1050
rect 25510 1030 25520 1050
rect 25330 1020 25520 1030
rect 27020 -425 27125 1100
rect 27020 -445 27245 -425
rect 26820 -1800 26865 -1790
rect 26820 -1820 26830 -1800
rect 26855 -1820 26865 -1800
rect 26820 -1830 26865 -1820
rect 17955 -2040 18005 -2025
rect 17955 -2060 17970 -2040
rect 17990 -2060 18005 -2040
rect 17955 -2075 18005 -2060
rect -85 -2125 -35 -2110
rect -85 -2145 -70 -2125
rect -50 -2145 -35 -2125
rect 17875 -2130 18105 -2095
rect -85 -2440 -35 -2145
rect 17955 -2165 18005 -2150
rect 17955 -2185 17970 -2165
rect 17990 -2185 18005 -2165
rect -85 -2480 50 -2440
rect 17955 -2480 18005 -2185
rect 17955 -2520 18090 -2480
rect 17615 -2560 17655 -2545
rect 17615 -2580 17625 -2560
rect 17645 -2580 17655 -2560
rect 17615 -2590 17655 -2580
rect 17920 -2555 17965 -2545
rect 17920 -2580 17930 -2555
rect 17955 -2580 17965 -2555
rect 17920 -2590 17965 -2580
rect 17615 -2765 17970 -2755
rect 17615 -2795 17625 -2765
rect 17665 -2770 17970 -2765
rect 17665 -2790 17930 -2770
rect 17950 -2790 17970 -2770
rect 17665 -2795 17970 -2790
rect 17615 -2805 17970 -2795
rect 8985 -3920 9090 -3900
rect 8985 -3990 9005 -3920
rect 9070 -3990 9090 -3920
rect 8985 -4300 9090 -3990
rect 7365 -4340 9090 -4300
rect 27020 -3960 27125 -3940
rect 27020 -4030 27040 -3960
rect 27105 -4030 27125 -3960
rect 27020 -4340 27125 -4030
rect 25405 -4380 27125 -4340
<< viali >>
rect 8790 1485 8815 1505
rect 9000 1215 9065 1285
rect 7450 1080 7470 1100
rect 17560 -1350 17600 -1310
rect 8610 -1455 8630 -1435
rect 9150 -1455 9170 -1435
rect 8795 -1780 8820 -1760
rect 26830 1445 26855 1465
rect 27040 1175 27105 1245
rect 25490 1030 25510 1050
rect 26830 -1820 26855 -1800
rect 17625 -2580 17645 -2560
rect 17930 -2580 17955 -2555
rect 17625 -2795 17665 -2765
rect 17930 -2790 17950 -2770
rect 9005 -3990 9070 -3920
rect 27040 -4030 27105 -3960
<< metal1 >>
rect 4610 5375 22855 5560
rect -235 3285 35 3325
rect 4610 3305 4710 5375
rect -235 -2785 -200 3285
rect 4610 3250 5620 3305
rect 4610 3075 4710 3250
rect 5520 3075 5620 3250
rect 8780 1510 8830 1515
rect 8780 1480 8785 1510
rect 8820 1480 8830 1510
rect 8780 1455 8830 1480
rect 7440 1435 8830 1455
rect 7440 1110 7460 1435
rect 7440 1100 7480 1110
rect 7240 1070 7290 1090
rect 7440 1080 7450 1100
rect 7470 1080 7480 1100
rect 7440 1070 7480 1080
rect 6220 205 6770 930
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 6220 110 6770 120
rect -120 -5 25 15
rect -120 -2155 -75 -5
rect 6220 -90 6770 -80
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -970 6770 -175
rect 5335 -1505 6770 -970
rect 7365 -1425 7385 25
rect 8780 -100 8830 1435
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 13560 1060 13660 5375
rect 22645 3320 22855 5375
rect 13560 865 13570 1060
rect 13650 865 13660 1060
rect 13560 580 13660 865
rect 17805 3245 18075 3285
rect 8780 -135 10025 -100
rect 7365 -1435 8640 -1425
rect 7365 -1445 8610 -1435
rect 8600 -1455 8610 -1445
rect 8630 -1455 8640 -1435
rect 8600 -1465 8640 -1455
rect 5335 -1975 5645 -1505
rect 8780 -1755 8830 -135
rect 17550 -1310 17610 -1300
rect 17550 -1350 17560 -1310
rect 17600 -1350 17610 -1310
rect 17550 -1360 17610 -1350
rect 9140 -1435 12755 -1425
rect 9140 -1455 9150 -1435
rect 9170 -1445 12755 -1435
rect 9170 -1455 9180 -1445
rect 9140 -1465 9180 -1455
rect 8780 -1785 8790 -1755
rect 8825 -1785 8830 -1755
rect 8780 -1790 8830 -1785
rect 8785 -1885 8830 -1825
rect -120 -2195 45 -2155
rect 4625 -2285 5645 -1975
rect 12720 -2120 12755 -1445
rect 12720 -2160 17655 -2120
rect 4625 -2405 4725 -2285
rect 5545 -2405 5645 -2285
rect 17615 -2560 17655 -2160
rect 17615 -2580 17625 -2560
rect 17645 -2580 17655 -2560
rect 17615 -2590 17655 -2580
rect 17615 -2765 17675 -2755
rect -235 -2820 25 -2785
rect 17615 -2795 17625 -2765
rect 17665 -2795 17675 -2765
rect 17615 -2805 17675 -2795
rect 17805 -2825 17840 3245
rect 22645 3215 23660 3320
rect 22645 3030 22780 3215
rect 23525 3035 23660 3215
rect 26820 1470 26865 1475
rect 26820 1440 26825 1470
rect 26860 1440 26865 1470
rect 26820 1415 26865 1440
rect 25480 1395 26865 1415
rect 25480 1060 25500 1395
rect 25480 1050 25520 1060
rect 25280 1030 25330 1050
rect 25480 1030 25490 1050
rect 25510 1030 25520 1050
rect 25480 1020 25520 1030
rect 24260 165 24810 890
rect 24260 80 24270 165
rect 24800 80 24810 165
rect 24260 70 24810 80
rect 17920 -45 18065 -25
rect 17920 -2195 17965 -45
rect 24260 -130 24810 -120
rect 24260 -215 24270 -130
rect 24800 -215 24810 -130
rect 24260 -1010 24810 -215
rect 23375 -1545 24810 -1010
rect 26820 -140 26865 1395
rect 27030 1245 27115 1255
rect 27030 1175 27040 1245
rect 27105 1175 27115 1245
rect 27030 1165 27115 1175
rect 26820 -175 27245 -140
rect 23375 -2015 23685 -1545
rect 26820 -1795 26865 -175
rect 26820 -1825 26825 -1795
rect 26860 -1825 26865 -1795
rect 26820 -1830 26865 -1825
rect 26820 -1925 26865 -1865
rect 17920 -2235 18085 -2195
rect 17920 -2555 17965 -2235
rect 22665 -2325 23685 -2015
rect 22665 -2445 22765 -2325
rect 23585 -2445 23685 -2325
rect 17920 -2580 17930 -2555
rect 17955 -2580 17965 -2555
rect 17920 -2590 17965 -2580
rect 17915 -2765 17970 -2755
rect 17915 -2795 17925 -2765
rect 17955 -2795 17970 -2765
rect 17915 -2805 17970 -2795
rect 17805 -2860 18065 -2825
rect 8995 -3920 9080 -3910
rect 8995 -3990 9005 -3920
rect 9070 -3990 9080 -3920
rect 8995 -4000 9080 -3990
rect 27030 -3960 27115 -3950
rect 27030 -4030 27040 -3960
rect 27105 -4030 27115 -3960
rect 27030 -4040 27115 -4030
rect 7405 -5485 18080 -5465
<< via1 >>
rect 8785 1505 8820 1510
rect 8785 1485 8790 1505
rect 8790 1485 8815 1505
rect 8815 1485 8820 1505
rect 8785 1480 8820 1485
rect 6230 120 6760 205
rect 6230 -175 6760 -90
rect 9000 1215 9065 1285
rect 13570 865 13650 1060
rect 17560 -1350 17600 -1310
rect 8790 -1760 8825 -1755
rect 8790 -1780 8795 -1760
rect 8795 -1780 8820 -1760
rect 8820 -1780 8825 -1760
rect 8790 -1785 8825 -1780
rect 17625 -2795 17665 -2765
rect 26825 1465 26860 1470
rect 26825 1445 26830 1465
rect 26830 1445 26855 1465
rect 26855 1445 26860 1465
rect 26825 1440 26860 1445
rect 24270 80 24800 165
rect 24270 -215 24800 -130
rect 27040 1175 27105 1245
rect 26825 -1800 26860 -1795
rect 26825 -1820 26830 -1800
rect 26830 -1820 26855 -1800
rect 26855 -1820 26860 -1800
rect 26825 -1825 26860 -1820
rect 17925 -2770 17955 -2765
rect 17925 -2790 17930 -2770
rect 17930 -2790 17950 -2770
rect 17950 -2790 17955 -2770
rect 17925 -2795 17955 -2790
rect 9005 -3990 9070 -3920
rect 27040 -4030 27105 -3960
<< metal2 >>
rect 4005 5355 22585 5560
rect 4005 3075 4540 5355
rect -235 2720 15 2760
rect -235 -3350 -200 2720
rect 8780 1510 8825 1515
rect 8780 1480 8785 1510
rect 8820 1480 8825 1510
rect 8780 1475 8825 1480
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 4005 685 4425 835
rect 4005 470 4270 685
rect 12960 585 13395 5355
rect 22045 3035 22585 5355
rect 17805 2680 18055 2720
rect 13560 1060 13660 1070
rect 13560 865 13570 1060
rect 13650 865 13660 1060
rect 13560 855 13660 865
rect 4005 405 4015 470
rect 4260 405 4270 470
rect 4005 395 4270 405
rect 6220 205 6770 215
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 6220 110 6770 120
rect -120 -5 25 15
rect -120 -2720 -75 -5
rect 4025 -65 4355 -55
rect 4025 -145 4035 -65
rect 4345 -145 4355 -65
rect 4025 -2405 4355 -145
rect 6220 -90 6770 -80
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -185 6770 -175
rect 7365 -1425 7385 25
rect 17550 -1310 17610 -1300
rect 17550 -1350 17560 -1310
rect 17600 -1350 17610 -1310
rect 17550 -1360 17610 -1350
rect 7365 -1445 12755 -1425
rect 8785 -1755 8830 -1750
rect 8785 -1785 8790 -1755
rect 8825 -1785 8830 -1755
rect 8785 -1790 8830 -1785
rect 12720 -2120 12755 -1445
rect 12720 -2160 17655 -2120
rect -120 -2760 30 -2720
rect 17615 -2755 17655 -2160
rect 17615 -2765 17675 -2755
rect 17615 -2795 17625 -2765
rect 17665 -2795 17675 -2765
rect 17615 -2805 17675 -2795
rect -235 -3390 60 -3350
rect 17805 -3390 17840 2680
rect 26820 1470 26865 1475
rect 26820 1440 26825 1470
rect 26860 1440 26865 1470
rect 26820 1435 26865 1440
rect 27030 1245 27115 1255
rect 27030 1175 27040 1245
rect 27105 1175 27115 1245
rect 27030 1165 27115 1175
rect 22045 645 22465 795
rect 22045 430 22310 645
rect 22045 365 22055 430
rect 22300 365 22310 430
rect 22045 355 22310 365
rect 24260 165 24810 175
rect 24260 80 24270 165
rect 24800 80 24810 165
rect 24260 70 24810 80
rect 17920 -45 18065 -25
rect 17920 -2755 17965 -45
rect 22065 -105 22395 -95
rect 22065 -185 22075 -105
rect 22385 -185 22395 -105
rect 22065 -2445 22395 -185
rect 24260 -130 24810 -120
rect 24260 -215 24270 -130
rect 24800 -215 24810 -130
rect 24260 -225 24810 -215
rect 26820 -1795 26865 -1790
rect 26820 -1825 26825 -1795
rect 26860 -1825 26865 -1795
rect 26820 -1830 26865 -1825
rect 17915 -2760 17970 -2755
rect 17915 -2765 18070 -2760
rect 17915 -2795 17925 -2765
rect 17955 -2795 18070 -2765
rect 17915 -2800 18070 -2795
rect 17915 -2805 17970 -2800
rect 17805 -3430 18100 -3390
rect 8995 -3920 9080 -3910
rect 8995 -3990 9005 -3920
rect 9070 -3990 9080 -3920
rect 8995 -4000 9080 -3990
rect 27030 -3960 27115 -3950
rect 27030 -4030 27040 -3960
rect 27105 -4030 27115 -3960
rect 27030 -4040 27115 -4030
rect 7405 -5485 18080 -5465
<< via2 >>
rect 8785 1480 8820 1510
rect 9000 1215 9065 1285
rect 13570 865 13650 1060
rect 4015 405 4260 470
rect 6230 120 6760 205
rect 4035 -145 4345 -65
rect 6230 -175 6760 -90
rect 17560 -1350 17600 -1310
rect 8790 -1785 8825 -1755
rect 26825 1440 26860 1470
rect 27040 1175 27105 1245
rect 22055 365 22300 430
rect 24270 80 24800 165
rect 22075 -185 22385 -105
rect 24270 -215 24800 -130
rect 26825 -1825 26860 -1795
rect 9005 -3990 9070 -3920
rect 27040 -4030 27105 -3960
<< metal3 >>
rect -250 3155 1405 3210
rect -250 -2270 -190 3155
rect 17790 3115 19445 3170
rect 8775 1510 8830 1585
rect 8775 1480 8785 1510
rect 8820 1480 8830 1510
rect 8775 1475 8830 1480
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 12445 1060 13660 1070
rect 12445 865 13570 1060
rect 13650 865 13660 1060
rect 12445 855 13660 865
rect 4005 470 4270 480
rect 4005 405 4015 470
rect 4260 405 4270 470
rect 4005 395 4270 405
rect 4025 -55 4270 395
rect 6220 205 6770 215
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 4025 -65 4355 -55
rect 4025 -145 4035 -65
rect 4345 -145 4355 -65
rect 4025 -155 4355 -145
rect 6220 -90 6770 120
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -185 6770 -175
rect 17790 -1300 17850 3115
rect 26815 1470 26870 1545
rect 26815 1440 26825 1470
rect 26860 1440 26870 1470
rect 26815 1435 26870 1440
rect 27030 1245 27115 1255
rect 27030 1175 27040 1245
rect 27105 1175 27115 1245
rect 27030 1165 27115 1175
rect 22045 430 22310 440
rect 22045 365 22055 430
rect 22300 365 22310 430
rect 22045 355 22310 365
rect 22065 -95 22310 355
rect 24260 165 24810 175
rect 24260 80 24270 165
rect 24800 80 24810 165
rect 22065 -105 22395 -95
rect 22065 -185 22075 -105
rect 22385 -185 22395 -105
rect 22065 -195 22395 -185
rect 24260 -130 24810 80
rect 24260 -215 24270 -130
rect 24800 -215 24810 -130
rect 24260 -225 24810 -215
rect 17550 -1310 17850 -1300
rect 17550 -1350 17560 -1310
rect 17600 -1350 17850 -1310
rect 17550 -1360 17850 -1350
rect 8780 -1755 8835 -1750
rect 8780 -1785 8790 -1755
rect 8825 -1785 8835 -1755
rect 8780 -1855 8835 -1785
rect -255 -2320 1260 -2270
rect 17790 -2310 17850 -1360
rect 26815 -1795 26870 -1790
rect 26815 -1825 26825 -1795
rect 26860 -1825 26870 -1795
rect 26815 -1895 26870 -1825
rect 17790 -2360 19300 -2310
rect 8995 -3920 9080 -3910
rect 8995 -3990 9005 -3920
rect 9070 -3990 9080 -3920
rect 8995 -4000 9080 -3990
rect 27030 -3960 27115 -3950
rect 27030 -4030 27040 -3960
rect 27105 -4030 27115 -3960
rect 27030 -4040 27115 -4030
<< via3 >>
rect 9000 1215 9065 1285
rect 27040 1175 27105 1245
rect 9005 -3990 9070 -3920
rect 27040 -4030 27105 -3960
<< metal4 >>
rect 8980 1285 9085 1840
rect 8980 1215 9000 1285
rect 9065 1215 9085 1285
rect 8980 -1580 9085 1215
rect 27020 1245 27125 1800
rect 27020 1175 27040 1245
rect 27105 1175 27125 1245
rect 8985 -2125 9090 -1580
rect 27020 -2165 27125 1175
rect 8985 -3920 9090 -3320
rect 8985 -3990 9005 -3920
rect 9070 -3990 9090 -3920
rect 8985 -4065 9090 -3990
rect 27020 -3960 27125 -3360
rect 27020 -4030 27040 -3960
rect 27105 -4030 27125 -3960
rect 27020 -4105 27125 -4030
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_1
timestamp 1620752477
transform 1 0 3950 0 1 -4910
box -3935 -575 4700 4735
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_3
timestamp 1620752477
transform 1 0 21990 0 1 -4950
box -3935 -575 4700 4735
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_0
timestamp 1620752477
transform 1 0 3930 0 1 570
box -3935 -575 4700 4735
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_2
timestamp 1620752477
transform 1 0 21970 0 1 530
box -3935 -575 4700 4735
use middle_ping_pong_amplifier  middle_ping_pong_amplifier_0
timestamp 1620752477
transform 1 0 12905 0 1 -1890
box -3700 -30 4680 3175
use cap8to1  cap8to1_3
timestamp 1620749136
transform 1 0 26800 0 1 1455
box 5 30 3785 1860
use cap8to1  cap8to1_1
timestamp 1620749136
transform 1 0 8760 0 1 1495
box 5 30 3785 1860
use cap8to1  cap8to1_0
timestamp 1620749136
transform 1 0 8765 0 1 -3670
box 5 30 3785 1860
use cap8to1  cap8to1_2
timestamp 1620749136
transform 1 0 26805 0 1 -3710
box 5 30 3785 1860
<< end >>
