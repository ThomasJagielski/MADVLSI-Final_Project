**.subckt counter-bn_lvs
X16 Qn8 __UNCONNECTED_PIN__0 net1 net2 P C dff
X17 net1 Qn8 __UNCONNECTED_PIN__1 Q7 C P dff
X20 Q7 net2 VDD GND inverter
X24 net1 Q8 VDD GND inverter
**.ends

* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/dff.sym # of pins=6

.subckt dff  D Qn Q CLK Preset Clear
*.ipin D
*.iopin CLK
*.opin Qn
*.opin Q
*.ipin Preset
*.ipin Clear
X6 D CLK net4 VDD GND nand2
X7 net1 CLK net2 VDD GND nand2
X8 Q net3 Qn VDD GND nand2
X9 net5 Qn Q VDD GND nand2
X10 D net1 VDD GND inverter
X1 VDD Preset GND net5 net4 and2
X2 VDD net2 GND net3 Clear and2
.ends


* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/inverter.sym # of
*+ pins=4

.subckt inverter  A Y VP VN
*.ipin A
*.iopin VP
*.iopin VN
*.opin Y
XM1 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 Y A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/nand2.sym # of pins=5

.subckt nand2  A B Y VP VN
*.ipin A
*.opin Y
*.ipin B
*.iopin VP
*.iopin VP
*.iopin VN
*.iopin VN
XM1 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 VP B Y VP sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 B Y VN sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net1 A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/and2.sym # of pins=5

.subckt and2  VP A VN Y B
*.iopin VP
*.iopin VN
*.ipin A
*.ipin B
*.opin Y
X1 A B net1 VP VN nand2
X2 net1 Y VP VN inverter
.ends

.GLOBAL VDD
.GLOBAL GND
** flattened .save nodes
.end
