* NGSPICE file created from decimation_filter.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt decimation_filter DATA[0] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15]
+ DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] data_en
+ dec_rate[0] dec_rate[10] dec_rate[11] dec_rate[12] dec_rate[13] dec_rate[14] dec_rate[15]
+ dec_rate[1] dec_rate[2] dec_rate[3] dec_rate[4] dec_rate[5] dec_rate[6] dec_rate[7]
+ dec_rate[8] dec_rate[9] mclk1 mdata1 reset VPWR VGND
X_3155_ _4153_/A VGND VGND VPWR VPWR _3660_/A sky130_fd_sc_hd__clkbuf_2
X_3086_ _3086_/A VGND VGND VPWR VPWR _3086_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3988_ _3831_/A _3994_/B _3994_/A _3827_/A VGND VGND VPWR VPWR _3989_/B sky130_fd_sc_hd__a31o_1
XFILLER_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2939_ _2939_/A VGND VGND VPWR VPWR _3158_/B sky130_fd_sc_hd__inv_2
X_4609_ _4621_/A VGND VGND VPWR VPWR _4614_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer7 _3351_/B VGND VGND VPWR VPWR _3388_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4960_ _5018_/CLK _4960_/D VGND VGND VPWR VPWR _4960_/Q sky130_fd_sc_hd__dfxtp_1
X_4891_ _5047_/CLK _4891_/D VGND VGND VPWR VPWR _4891_/Q sky130_fd_sc_hd__dfxtp_1
X_3911_ _3911_/A VGND VGND VPWR VPWR _3913_/A sky130_fd_sc_hd__inv_2
XFILLER_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3842_ _3842_/A VGND VGND VPWR VPWR _4000_/A sky130_fd_sc_hd__inv_2
X_3773_ _3604_/B _5035_/Q _3604_/B _5035_/Q VGND VGND VPWR VPWR _3923_/B sky130_fd_sc_hd__a2bb2o_1
X_2724_ _2801_/A _2722_/X _2723_/X VGND VGND VPWR VPWR _2735_/A sky130_fd_sc_hd__o21a_1
X_2655_ _2691_/A _2624_/B _2590_/D VGND VGND VPWR VPWR _2656_/D sky130_fd_sc_hd__o21a_1
X_4325_ _4325_/A VGND VGND VPWR VPWR _4326_/A sky130_fd_sc_hd__buf_1
X_2586_ _2775_/A VGND VGND VPWR VPWR _2590_/C sky130_fd_sc_hd__clkbuf_2
X_4256_ _3728_/B _4980_/Q _4255_/Y VGND VGND VPWR VPWR _4257_/A sky130_fd_sc_hd__o21ai_1
X_4187_ _4192_/A _4192_/B VGND VGND VPWR VPWR _4193_/B sky130_fd_sc_hd__or2_1
X_3207_ _3212_/A _3207_/B VGND VGND VPWR VPWR _3207_/X sky130_fd_sc_hd__or2_1
X_3138_ _5132_/Q VGND VGND VPWR VPWR _3138_/Y sky130_fd_sc_hd__inv_2
X_3069_ _3327_/A _4721_/B VGND VGND VPWR VPWR _3069_/Y sky130_fd_sc_hd__nor2_2
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2440_ _4664_/A _2440_/B VGND VGND VPWR VPWR _2440_/X sky130_fd_sc_hd__or2_1
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4110_ _4101_/Y _4271_/A _4266_/A _4109_/X VGND VGND VPWR VPWR _4253_/A sky130_fd_sc_hd__o31a_1
X_5090_ _3391_/X _5090_/D VGND VGND VPWR VPWR _5090_/Q sky130_fd_sc_hd__dfxtp_2
X_4041_ _4041_/A _4041_/B VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__or2_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4943_ _5018_/CLK _4943_/D VGND VGND VPWR VPWR _4943_/Q sky130_fd_sc_hd__dfxtp_1
X_4874_ _5028_/CLK _4874_/D VGND VGND VPWR VPWR _4874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3825_ _3825_/A _5015_/Q VGND VGND VPWR VPWR _3825_/Y sky130_fd_sc_hd__nor2_4
X_3756_ _5040_/Q VGND VGND VPWR VPWR _3756_/Y sky130_fd_sc_hd__inv_2
X_2707_ _2772_/A VGND VGND VPWR VPWR _2707_/X sky130_fd_sc_hd__buf_1
X_3687_ _3692_/A _3687_/B VGND VGND VPWR VPWR _4998_/D sky130_fd_sc_hd__nor2_1
X_2638_ _2770_/A VGND VGND VPWR VPWR _2638_/X sky130_fd_sc_hd__clkbuf_2
X_2569_ _4958_/Q _4960_/Q _4959_/Q _4957_/Q VGND VGND VPWR VPWR _2603_/D sky130_fd_sc_hd__or4_4
X_4308_ _4814_/Q VGND VGND VPWR VPWR _4458_/A sky130_fd_sc_hd__inv_2
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4239_ _4250_/A _4084_/B _4116_/Y VGND VGND VPWR VPWR _4240_/B sky130_fd_sc_hd__o21ai_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3610_ _4921_/Q VGND VGND VPWR VPWR _3611_/B sky130_fd_sc_hd__inv_2
X_4590_ _4398_/Y _4588_/Y _4406_/A _3996_/X _4589_/Y VGND VGND VPWR VPWR _4868_/D
+ sky130_fd_sc_hd__o311a_1
X_3541_ _3481_/A _3540_/Y _5056_/Q _3540_/Y VGND VGND VPWR VPWR _3542_/D sky130_fd_sc_hd__a2bb2o_1
X_3472_ _5060_/Q VGND VGND VPWR VPWR _3486_/A sky130_fd_sc_hd__inv_2
X_2423_ _4575_/A VGND VGND VPWR VPWR _2423_/X sky130_fd_sc_hd__buf_2
X_5073_ _3442_/X _5073_/D VGND VGND VPWR VPWR _5073_/Q sky130_fd_sc_hd__dfxtp_1
X_4024_ _4024_/A VGND VGND VPWR VPWR _4025_/B sky130_fd_sc_hd__inv_2
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4926_ _5047_/CLK _4926_/D VGND VGND VPWR VPWR _4926_/Q sky130_fd_sc_hd__dfxtp_1
X_4857_ _5047_/CLK _4857_/D VGND VGND VPWR VPWR _4857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3808_ _3808_/A _3967_/A VGND VGND VPWR VPWR _3809_/B sky130_fd_sc_hd__or2_1
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4788_ _2563_/X _4788_/D VGND VGND VPWR VPWR _4788_/Q sky130_fd_sc_hd__dfxtp_1
X_3739_ _4864_/Q VGND VGND VPWR VPWR _3740_/B sky130_fd_sc_hd__inv_2
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2972_ _2972_/A VGND VGND VPWR VPWR _2972_/X sky130_fd_sc_hd__clkbuf_2
X_4711_ _4711_/A VGND VGND VPWR VPWR _4714_/A sky130_fd_sc_hd__inv_2
X_4642_ _4644_/A _4722_/A VGND VGND VPWR VPWR _4830_/D sky130_fd_sc_hd__nor2_1
X_4573_ _4637_/B _4834_/Q _4578_/B VGND VGND VPWR VPWR _4574_/A sky130_fd_sc_hd__o21ai_1
X_3524_ _3523_/A _3523_/B _3523_/Y VGND VGND VPWR VPWR _3525_/B sky130_fd_sc_hd__a21oi_1
X_3455_ _3455_/A VGND VGND VPWR VPWR _3455_/X sky130_fd_sc_hd__buf_1
X_2406_ _2406_/A VGND VGND VPWR VPWR _2406_/Y sky130_fd_sc_hd__inv_2
X_3386_ _3396_/A VGND VGND VPWR VPWR _3386_/X sky130_fd_sc_hd__buf_1
XFILLER_69_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5125_ _3211_/X _5125_/D VGND VGND VPWR VPWR _5125_/Q sky130_fd_sc_hd__dfxtp_1
X_5056_ _5063_/CLK _5056_/D VGND VGND VPWR VPWR _5056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4007_ _4900_/Q _3837_/Y _3659_/B _5011_/Q VGND VGND VPWR VPWR _4008_/B sky130_fd_sc_hd__o22a_1
XFILLER_55_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4909_ _5028_/CLK _4909_/D VGND VGND VPWR VPWR _4909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 _4596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3240_ _3235_/A _3235_/B _3223_/X _3235_/Y VGND VGND VPWR VPWR _5119_/D sky130_fd_sc_hd__o211a_1
XFILLER_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3171_ _2942_/Y _3170_/Y _2942_/A _3170_/A _3660_/A VGND VGND VPWR VPWR _5134_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer17 _3341_/B VGND VGND VPWR VPWR _3414_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer39 _3347_/B VGND VGND VPWR VPWR _3395_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer28 _3355_/B VGND VGND VPWR VPWR _3376_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2955_ _5093_/Q _2952_/X _3351_/A _2954_/Y VGND VGND VPWR VPWR _2956_/A sky130_fd_sc_hd__o22a_1
X_2886_ _5054_/Q _2885_/A _3479_/A _2885_/Y VGND VGND VPWR VPWR _2886_/X sky130_fd_sc_hd__a22o_1
X_4625_ _4626_/A _4625_/B VGND VGND VPWR VPWR _4844_/D sky130_fd_sc_hd__nor2_1
X_4556_ _4552_/A _4552_/B _4526_/X _4552_/Y VGND VGND VPWR VPWR _4877_/D sky130_fd_sc_hd__o211a_1
X_3507_ _3508_/A _3507_/B VGND VGND VPWR VPWR _3507_/Y sky130_fd_sc_hd__nor2_1
X_4487_ _4578_/A _4487_/B _4487_/C VGND VGND VPWR VPWR _4895_/D sky130_fd_sc_hd__and3_1
X_3438_ _3333_/A _3438_/A2 _3431_/X _3434_/Y VGND VGND VPWR VPWR _5075_/D sky130_fd_sc_hd__a211oi_1
X_3369_ _3382_/A VGND VGND VPWR VPWR _3369_/X sky130_fd_sc_hd__buf_1
X_5108_ _3289_/X _5108_/D VGND VGND VPWR VPWR _5108_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5039_ _5047_/CLK _5039_/D VGND VGND VPWR VPWR _5039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput20 _4782_/Q VGND VGND VPWR VPWR DATA[10] sky130_fd_sc_hd__clkbuf_2
Xoutput31 _4778_/Q VGND VGND VPWR VPWR DATA[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2740_ _2643_/A _2709_/X _2710_/X VGND VGND VPWR VPWR _2742_/C sky130_fd_sc_hd__o21a_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2671_ _4941_/Q _2630_/B _2590_/C VGND VGND VPWR VPWR _2674_/C sky130_fd_sc_hd__o21a_1
X_4410_ _4410_/A VGND VGND VPWR VPWR _4410_/Y sky130_fd_sc_hd__inv_2
X_4341_ _4348_/A _4844_/Q _4348_/A _4844_/Q VGND VGND VPWR VPWR _4534_/A sky130_fd_sc_hd__a2bb2o_1
X_4272_ _4108_/A _4271_/Y _4264_/X _4266_/X VGND VGND VPWR VPWR _4902_/D sky130_fd_sc_hd__o211a_1
X_3223_ _3375_/A VGND VGND VPWR VPWR _3223_/X sky130_fd_sc_hd__clkbuf_2
X_3154_ _4500_/A VGND VGND VPWR VPWR _4153_/A sky130_fd_sc_hd__clkbuf_2
X_3085_ _5103_/Q VGND VGND VPWR VPWR _3086_/A sky130_fd_sc_hd__inv_2
XFILLER_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3987_ _3987_/A VGND VGND VPWR VPWR _3994_/A sky130_fd_sc_hd__inv_2
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2938_ _3356_/A _2937_/X _5098_/Q _5135_/Q VGND VGND VPWR VPWR _2939_/A sky130_fd_sc_hd__o22a_1
X_2869_ _5057_/Q VGND VGND VPWR VPWR _3483_/A sky130_fd_sc_hd__clkbuf_2
X_4608_ _4608_/A _4608_/B VGND VGND VPWR VPWR _4858_/D sky130_fd_sc_hd__nor2_1
X_4539_ _4575_/A VGND VGND VPWR VPWR _4539_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer8 _3351_/B VGND VGND VPWR VPWR _3383_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3910_ _3909_/Y _3897_/A _3462_/X _3905_/X VGND VGND VPWR VPWR _4965_/D sky130_fd_sc_hd__o211a_1
X_4890_ _5047_/CLK _4890_/D VGND VGND VPWR VPWR _4890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3841_ _3656_/B _5012_/Q _3840_/Y VGND VGND VPWR VPWR _3842_/A sky130_fd_sc_hd__o21ai_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3772_ _3772_/A VGND VGND VPWR VPWR _3774_/A sky130_fd_sc_hd__inv_2
X_2723_ _2788_/A VGND VGND VPWR VPWR _2723_/X sky130_fd_sc_hd__buf_1
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2654_ _4949_/Q VGND VGND VPWR VPWR _2691_/A sky130_fd_sc_hd__clkbuf_2
X_2585_ _2585_/A VGND VGND VPWR VPWR _2775_/A sky130_fd_sc_hd__inv_2
X_4324_ _4810_/Q VGND VGND VPWR VPWR _4325_/A sky130_fd_sc_hd__inv_2
X_4255_ _4255_/A _4255_/B VGND VGND VPWR VPWR _4255_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4186_ _4181_/A _4181_/B _4177_/X _4181_/Y VGND VGND VPWR VPWR _4926_/D sky130_fd_sc_hd__o211a_1
X_3206_ _3222_/A VGND VGND VPWR VPWR _3206_/X sky130_fd_sc_hd__buf_1
X_3137_ _5095_/Q VGND VGND VPWR VPWR _3353_/A sky130_fd_sc_hd__clkinv_1
XFILLER_67_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3068_ _5106_/Q VGND VGND VPWR VPWR _4721_/B sky130_fd_sc_hd__inv_2
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4040_ _4040_/A _4192_/B VGND VGND VPWR VPWR _4041_/B sky130_fd_sc_hd__or2_1
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4942_ _5018_/CLK _4942_/D VGND VGND VPWR VPWR _4942_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4873_ _5028_/CLK _4873_/D VGND VGND VPWR VPWR _4873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3824_ _3824_/A _5016_/Q VGND VGND VPWR VPWR _3824_/Y sky130_fd_sc_hd__nor2_1
X_3755_ _3595_/B _5039_/Q _3595_/B _5039_/Q VGND VGND VPWR VPWR _3909_/A sky130_fd_sc_hd__a2bb2o_1
X_3686_ _4887_/Q VGND VGND VPWR VPWR _3687_/B sky130_fd_sc_hd__inv_2
X_2706_ _2666_/A _2705_/X _2693_/X VGND VGND VPWR VPWR _2715_/A sky130_fd_sc_hd__o21a_1
X_2637_ _4942_/Q _2637_/B _2637_/C _2637_/D VGND VGND VPWR VPWR _2770_/A sky130_fd_sc_hd__nor4_2
X_2568_ _4956_/Q _4955_/Q _2567_/X VGND VGND VPWR VPWR _2573_/B sky130_fd_sc_hd__or3b_1
X_4307_ _4455_/A _4853_/Q _4455_/A _4853_/Q VGND VGND VPWR VPWR _4510_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2499_ _2498_/Y _4754_/A _2486_/X _2492_/X VGND VGND VPWR VPWR _4804_/D sky130_fd_sc_hd__o211a_1
X_4238_ _4238_/A VGND VGND VPWR VPWR _4240_/A sky130_fd_sc_hd__inv_2
X_4169_ _4031_/B _4168_/Y _4030_/A _4168_/A _4151_/X VGND VGND VPWR VPWR _4931_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ _2850_/A _3518_/X _3502_/Y VGND VGND VPWR VPWR _3540_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3471_ _3320_/X _3471_/A2 _5064_/Q _3471_/B2 _3359_/X VGND VGND VPWR VPWR _5064_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2422_ _2422_/A VGND VGND VPWR VPWR _2422_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5072_ _3445_/X _5072_/D VGND VGND VPWR VPWR _5072_/Q sky130_fd_sc_hd__dfxtp_1
X_4023_ _3675_/B _5003_/Q _4892_/Q _4022_/Y VGND VGND VPWR VPWR _4024_/A sky130_fd_sc_hd__o22a_1
XFILLER_69_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4925_ _5047_/CLK _4925_/D VGND VGND VPWR VPWR _4925_/Q sky130_fd_sc_hd__dfxtp_1
X_4856_ _5047_/CLK _4856_/D VGND VGND VPWR VPWR _4856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3807_ _3632_/B _5023_/Q _3632_/B _5023_/Q VGND VGND VPWR VPWR _3967_/A sky130_fd_sc_hd__a2bb2o_1
X_4787_ _5018_/CLK _4787_/D VGND VGND VPWR VPWR _4787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3738_ _4621_/A VGND VGND VPWR VPWR _4601_/A sky130_fd_sc_hd__clkbuf_2
X_3669_ _3669_/A VGND VGND VPWR VPWR _3679_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2971_ _5127_/Q VGND VGND VPWR VPWR _2972_/A sky130_fd_sc_hd__inv_2
X_4710_ _4636_/B _3049_/Y _4379_/X _5110_/Q VGND VGND VPWR VPWR _4711_/A sky130_fd_sc_hd__o22a_1
X_4641_ _4644_/A _4721_/A VGND VGND VPWR VPWR _4831_/D sky130_fd_sc_hd__nor2_1
X_4572_ _4577_/A _4577_/B VGND VGND VPWR VPWR _4578_/B sky130_fd_sc_hd__or2_1
X_3523_ _3523_/A _3523_/B VGND VGND VPWR VPWR _3523_/Y sky130_fd_sc_hd__nor2_1
X_3454_ _3327_/A _3454_/A2 _3431_/X _3451_/Y VGND VGND VPWR VPWR _5069_/D sky130_fd_sc_hd__a211oi_2
XFILLER_69_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2405_ _4652_/Y _4654_/Y _2416_/A _2404_/X VGND VGND VPWR VPWR _2406_/A sky130_fd_sc_hd__o31a_1
X_3385_ _3444_/A VGND VGND VPWR VPWR _3396_/A sky130_fd_sc_hd__buf_1
X_5124_ _3214_/X _5124_/D VGND VGND VPWR VPWR _5124_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5055_ _5063_/CLK _5055_/D VGND VGND VPWR VPWR _5055_/Q sky130_fd_sc_hd__dfxtp_1
X_4006_ _4900_/Q _3837_/Y _3839_/X _3996_/X _3840_/Y VGND VGND VPWR VPWR _4938_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4908_ _5028_/CLK _4908_/D VGND VGND VPWR VPWR _4908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4839_ _5028_/CLK _4839_/D VGND VGND VPWR VPWR _4839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 _4554_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3170_ _3170_/A VGND VGND VPWR VPWR _3170_/Y sky130_fd_sc_hd__inv_2
Xrebuffer18 _3353_/B VGND VGND VPWR VPWR _3381_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer29 _3339_/B VGND VGND VPWR VPWR _3423_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2954_ _5130_/Q VGND VGND VPWR VPWR _2954_/Y sky130_fd_sc_hd__inv_2
X_2885_ _2885_/A VGND VGND VPWR VPWR _2885_/Y sky130_fd_sc_hd__inv_2
X_4624_ _4626_/A _4624_/B VGND VGND VPWR VPWR _4845_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4555_ _4362_/A _4554_/Y _4359_/A _4554_/A _4539_/X VGND VGND VPWR VPWR _4878_/D
+ sky130_fd_sc_hd__o221a_1
X_3506_ input4/X VGND VGND VPWR VPWR _3506_/Y sky130_fd_sc_hd__inv_2
X_4486_ _4486_/A _4486_/B VGND VGND VPWR VPWR _4487_/C sky130_fd_sc_hd__nand2_1
X_3437_ _3442_/A VGND VGND VPWR VPWR _3437_/X sky130_fd_sc_hd__buf_1
X_3368_ _3368_/A VGND VGND VPWR VPWR _3382_/A sky130_fd_sc_hd__buf_1
X_5107_ _3297_/X _5107_/D VGND VGND VPWR VPWR _5107_/Q sky130_fd_sc_hd__dfxtp_1
X_3299_ _3312_/A VGND VGND VPWR VPWR _3299_/X sky130_fd_sc_hd__buf_1
X_5038_ _5047_/CLK _5038_/D VGND VGND VPWR VPWR _5038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput21 _4783_/Q VGND VGND VPWR VPWR DATA[11] sky130_fd_sc_hd__clkbuf_2
Xoutput32 _4779_/Q VGND VGND VPWR VPWR DATA[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2670_ _4938_/Q _2651_/X _2590_/B VGND VGND VPWR VPWR _2674_/B sky130_fd_sc_hd__o21a_1
X_4340_ _4806_/Q VGND VGND VPWR VPWR _4348_/A sky130_fd_sc_hd__inv_2
X_4271_ _4271_/A VGND VGND VPWR VPWR _4271_/Y sky130_fd_sc_hd__inv_2
X_3222_ _3222_/A VGND VGND VPWR VPWR _3222_/X sky130_fd_sc_hd__buf_1
X_3153_ _4176_/A VGND VGND VPWR VPWR _4500_/A sky130_fd_sc_hd__clkbuf_2
X_3084_ _5066_/Q VGND VGND VPWR VPWR _3324_/D sky130_fd_sc_hd__inv_1
XFILLER_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3986_ _3986_/A VGND VGND VPWR VPWR _3989_/A sky130_fd_sc_hd__inv_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2937_ _2937_/A VGND VGND VPWR VPWR _2937_/X sky130_fd_sc_hd__clkbuf_2
X_2868_ _5058_/Q _2867_/Y _5058_/Q _2867_/Y VGND VGND VPWR VPWR _2868_/X sky130_fd_sc_hd__o2bb2a_1
X_4607_ _4608_/A _4607_/B VGND VGND VPWR VPWR _4859_/D sky130_fd_sc_hd__nor2_1
X_2799_ _4965_/Q _2783_/X _2798_/X VGND VGND VPWR VPWR _2800_/D sky130_fd_sc_hd__o21a_1
X_4538_ _4538_/A VGND VGND VPWR VPWR _4538_/Y sky130_fd_sc_hd__inv_2
X_4469_ _4287_/Y _4486_/B _4486_/A _4468_/X VGND VGND VPWR VPWR _4480_/A sky130_fd_sc_hd__o31a_1
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer9 _3346_/B VGND VGND VPWR VPWR _3397_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3840_ _4900_/Q _3837_/Y _3839_/X VGND VGND VPWR VPWR _3840_/Y sky130_fd_sc_hd__o21ai_1
X_3771_ _3602_/B _5036_/Q _4925_/Q _3770_/Y VGND VGND VPWR VPWR _3772_/A sky130_fd_sc_hd__o22a_1
X_2722_ _2787_/A VGND VGND VPWR VPWR _2722_/X sky130_fd_sc_hd__buf_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2653_ _4940_/Q _2630_/B _2590_/C VGND VGND VPWR VPWR _2656_/C sky130_fd_sc_hd__o21a_1
X_2584_ _3517_/B _2584_/B _3517_/A VGND VGND VPWR VPWR _2585_/A sky130_fd_sc_hd__or3b_4
X_4323_ _4811_/Q VGND VGND VPWR VPWR _4619_/B sky130_fd_sc_hd__inv_2
X_4254_ _4097_/A _4260_/B _4260_/A _4093_/A VGND VGND VPWR VPWR _4255_/B sky130_fd_sc_hd__a31o_1
X_4185_ _4184_/A _4183_/Y _4184_/Y _4183_/A _4151_/X VGND VGND VPWR VPWR _4927_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3205_ _3199_/A _3199_/B _3186_/X _3199_/Y VGND VGND VPWR VPWR _5127_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3136_ _3349_/A _2968_/X _2985_/A _3134_/Y _3135_/X VGND VGND VPWR VPWR _3136_/X
+ sky130_fd_sc_hd__o221a_1
X_3067_ _5069_/Q VGND VGND VPWR VPWR _3327_/A sky130_fd_sc_hd__inv_2
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3969_ _3969_/A VGND VGND VPWR VPWR _3971_/A sky130_fd_sc_hd__inv_2
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4941_ _5018_/CLK _4941_/D VGND VGND VPWR VPWR _4941_/Q sky130_fd_sc_hd__dfxtp_1
X_4872_ _5028_/CLK _4872_/D VGND VGND VPWR VPWR _4872_/Q sky130_fd_sc_hd__dfxtp_1
X_3823_ _3645_/B _5017_/Q _3645_/B _5017_/Q VGND VGND VPWR VPWR _3986_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3754_ _3586_/B _5043_/Q _3586_/B _5043_/Q VGND VGND VPWR VPWR _3893_/B sky130_fd_sc_hd__a2bb2o_1
X_3685_ _3692_/A _3685_/B VGND VGND VPWR VPWR _4999_/D sky130_fd_sc_hd__nor2_1
X_2705_ _2770_/A VGND VGND VPWR VPWR _2705_/X sky130_fd_sc_hd__clkbuf_2
X_2636_ _2643_/A _2636_/B _4943_/Q _4944_/Q VGND VGND VPWR VPWR _2637_/C sky130_fd_sc_hd__or4_4
X_2567_ _4961_/Q VGND VGND VPWR VPWR _2567_/X sky130_fd_sc_hd__clkbuf_2
X_2498_ _4750_/X VGND VGND VPWR VPWR _2498_/Y sky130_fd_sc_hd__inv_2
X_4306_ _4815_/Q VGND VGND VPWR VPWR _4455_/A sky130_fd_sc_hd__inv_2
X_4237_ _4236_/Y _4224_/A _4220_/X _4232_/X VGND VGND VPWR VPWR _4912_/D sky130_fd_sc_hd__o211a_1
XFILLER_74_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4168_ _4168_/A VGND VGND VPWR VPWR _4168_/Y sky130_fd_sc_hd__inv_2
X_3119_ _3119_/A VGND VGND VPWR VPWR _3124_/A sky130_fd_sc_hd__inv_2
X_4099_ _4866_/Q _4099_/B VGND VGND VPWR VPWR _4099_/Y sky130_fd_sc_hd__nor2_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3470_ _4648_/A VGND VGND VPWR VPWR _3470_/X sky130_fd_sc_hd__buf_1
X_2421_ _4608_/B _2945_/X _2420_/X VGND VGND VPWR VPWR _2422_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5071_ _3448_/X _5071_/D VGND VGND VPWR VPWR _5071_/Q sky130_fd_sc_hd__dfxtp_1
X_4022_ _5003_/Q VGND VGND VPWR VPWR _4022_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4924_ _5047_/CLK _4924_/D VGND VGND VPWR VPWR _4924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4855_ _5047_/CLK _4855_/D VGND VGND VPWR VPWR _4855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4786_ _5047_/CLK _4786_/D VGND VGND VPWR VPWR _4786_/Q sky130_fd_sc_hd__dfxtp_1
X_3806_ _3806_/A VGND VGND VPWR VPWR _3808_/A sky130_fd_sc_hd__inv_2
X_3737_ _3737_/A VGND VGND VPWR VPWR _4621_/A sky130_fd_sc_hd__clkbuf_4
X_3668_ _3668_/A _3668_/B VGND VGND VPWR VPWR _5006_/D sky130_fd_sc_hd__nor2_1
X_3599_ _3599_/A _3599_/B VGND VGND VPWR VPWR _5037_/D sky130_fd_sc_hd__nor2_1
X_2619_ _4948_/Q _4952_/Q _4953_/Q VGND VGND VPWR VPWR _2620_/C sky130_fd_sc_hd__or3_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2970_ _5090_/Q VGND VGND VPWR VPWR _3348_/A sky130_fd_sc_hd__inv_6
X_4640_ _4644_/A _4640_/B VGND VGND VPWR VPWR _4832_/D sky130_fd_sc_hd__nor2_1
X_4571_ _4566_/A _4566_/B _4562_/X _4566_/Y VGND VGND VPWR VPWR _4873_/D sky130_fd_sc_hd__o211a_1
X_3522_ input9/X _3522_/B VGND VGND VPWR VPWR _3523_/B sky130_fd_sc_hd__or2_1
X_3453_ _3455_/A VGND VGND VPWR VPWR _3453_/X sky130_fd_sc_hd__buf_1
X_2404_ _4606_/B _2937_/X _4650_/Y _4605_/B _3147_/Y VGND VGND VPWR VPWR _2404_/X
+ sky130_fd_sc_hd__o32a_1
X_3384_ _3384_/A VGND VGND VPWR VPWR _3444_/A sky130_fd_sc_hd__buf_1
X_5123_ _3222_/X _5123_/D VGND VGND VPWR VPWR _5123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5054_ _5139_/CLK _5054_/D VGND VGND VPWR VPWR _5054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4005_ _3842_/A _4004_/Y _3978_/X _4000_/X VGND VGND VPWR VPWR _4939_/D sky130_fd_sc_hd__o211a_1
XFILLER_80_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4907_ _5018_/CLK _4907_/D VGND VGND VPWR VPWR _4907_/Q sky130_fd_sc_hd__dfxtp_1
X_4838_ _5028_/CLK _4838_/D VGND VGND VPWR VPWR _4838_/Q sky130_fd_sc_hd__dfxtp_1
X_4769_ _2830_/X _2821_/X _4770_/S VGND VGND VPWR VPWR _4786_/D sky130_fd_sc_hd__mux2_2
XFILLER_4_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 _4735_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer19 _3353_/B VGND VGND VPWR VPWR _3378_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_47_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2953_ _5093_/Q VGND VGND VPWR VPWR _3351_/A sky130_fd_sc_hd__clkinv_1
X_2884_ _5054_/Q VGND VGND VPWR VPWR _3479_/A sky130_fd_sc_hd__inv_2
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4623_ _4626_/A _4623_/B VGND VGND VPWR VPWR _4846_/D sky130_fd_sc_hd__nor2_1
X_4554_ _4554_/A VGND VGND VPWR VPWR _4554_/Y sky130_fd_sc_hd__inv_2
X_3505_ _3483_/A _3504_/X _5057_/Q _3504_/X VGND VGND VPWR VPWR _3544_/A sky130_fd_sc_hd__a2bb2o_1
X_4485_ _4287_/Y _4484_/Y _4287_/A _4484_/A _4269_/X VGND VGND VPWR VPWR _4896_/D
+ sky130_fd_sc_hd__o221a_1
X_3436_ _5076_/Q _3434_/Y _3435_/X _3436_/C1 VGND VGND VPWR VPWR _5076_/D sky130_fd_sc_hd__o211a_1
X_3367_ _5098_/Q _3366_/Y _3287_/X _3367_/C1 VGND VGND VPWR VPWR _5098_/D sky130_fd_sc_hd__o211a_1
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5106_ _3299_/X _5106_/D VGND VGND VPWR VPWR _5106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5037_ _5047_/CLK _5037_/D VGND VGND VPWR VPWR _5037_/Q sky130_fd_sc_hd__dfxtp_1
X_3298_ _3292_/A _3292_/B _3287_/X _3292_/Y VGND VGND VPWR VPWR _5107_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput22 _4784_/Q VGND VGND VPWR VPWR DATA[12] sky130_fd_sc_hd__clkbuf_2
Xoutput33 _4780_/Q VGND VGND VPWR VPWR DATA[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4270_ _4101_/Y _4268_/Y _4101_/A _4268_/A _4269_/X VGND VGND VPWR VPWR _4903_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_79_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3221_ _3129_/B _3220_/Y _3127_/A _3220_/A _3193_/X VGND VGND VPWR VPWR _5124_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_79_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3152_ _3370_/A VGND VGND VPWR VPWR _4176_/A sky130_fd_sc_hd__inv_2
X_3083_ _3083_/A VGND VGND VPWR VPWR _3083_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3985_ _3985_/A _3985_/B _3985_/C VGND VGND VPWR VPWR _4945_/D sky130_fd_sc_hd__and3_1
X_2936_ _5135_/Q VGND VGND VPWR VPWR _2937_/A sky130_fd_sc_hd__inv_2
X_2867_ _2864_/Y _3512_/B _3507_/B VGND VGND VPWR VPWR _2867_/Y sky130_fd_sc_hd__o21ai_1
X_4606_ _4608_/A _4606_/B VGND VGND VPWR VPWR _4860_/D sky130_fd_sc_hd__nor2_1
X_2798_ _2798_/A VGND VGND VPWR VPWR _2798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4537_ _4625_/B _4844_/Q _4536_/Y VGND VGND VPWR VPWR _4538_/A sky130_fd_sc_hd__o21ai_1
X_4468_ _4608_/B _4858_/Q _4285_/Y _4607_/B _4859_/Q VGND VGND VPWR VPWR _4468_/X
+ sky130_fd_sc_hd__o32a_1
X_3419_ _3426_/A VGND VGND VPWR VPWR _3419_/X sky130_fd_sc_hd__buf_1
X_4399_ _4721_/A _4831_/Q _4396_/Y _4398_/Y VGND VGND VPWR VPWR _4400_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3770_ _5036_/Q VGND VGND VPWR VPWR _3770_/Y sky130_fd_sc_hd__inv_2
X_2721_ _2721_/A _2756_/B VGND VGND VPWR VPWR _2721_/X sky130_fd_sc_hd__or2_1
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2652_ _4937_/Q _2651_/X _2590_/B VGND VGND VPWR VPWR _2656_/B sky130_fd_sc_hd__o21a_1
X_2583_ _2772_/A VGND VGND VPWR VPWR _2590_/B sky130_fd_sc_hd__clkbuf_2
X_4322_ _4811_/Q _4322_/B VGND VGND VPWR VPWR _4322_/Y sky130_fd_sc_hd__nor2_1
X_4253_ _4253_/A VGND VGND VPWR VPWR _4260_/A sky130_fd_sc_hd__inv_2
X_3204_ _3222_/A VGND VGND VPWR VPWR _3204_/X sky130_fd_sc_hd__buf_1
XFILLER_79_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4184_ _4184_/A VGND VGND VPWR VPWR _4184_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3135_ _3349_/A _2968_/X _3348_/A _2972_/X VGND VGND VPWR VPWR _3135_/X sky130_fd_sc_hd__a211o_1
X_3066_ _3292_/A VGND VGND VPWR VPWR _3103_/B sky130_fd_sc_hd__inv_2
XFILLER_23_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3968_ _3967_/Y _3956_/A _3939_/X _3963_/X VGND VGND VPWR VPWR _4949_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2919_ _3487_/A _2876_/X _2918_/X VGND VGND VPWR VPWR _2919_/Y sky130_fd_sc_hd__o21ai_1
X_3899_ _3899_/A _3899_/B VGND VGND VPWR VPWR _3899_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4940_ _5018_/CLK _4940_/D VGND VGND VPWR VPWR _4940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4871_ _5028_/CLK _4871_/D VGND VGND VPWR VPWR _4871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3822_ _3822_/A VGND VGND VPWR VPWR _3845_/A sky130_fd_sc_hd__inv_2
X_3753_ _3753_/A VGND VGND VPWR VPWR _3753_/Y sky130_fd_sc_hd__inv_2
X_3684_ _4888_/Q VGND VGND VPWR VPWR _3685_/B sky130_fd_sc_hd__inv_2
X_2704_ _2786_/A _2645_/X _2647_/X VGND VGND VPWR VPWR _2720_/A sky130_fd_sc_hd__o21a_1
X_2635_ _4946_/Q VGND VGND VPWR VPWR _2643_/A sky130_fd_sc_hd__clkbuf_2
X_4305_ _4305_/A _4305_/B VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__or2_1
X_2566_ _4950_/Q _4949_/Q VGND VGND VPWR VPWR _2632_/B sky130_fd_sc_hd__or2_2
X_2497_ _2497_/A VGND VGND VPWR VPWR _2497_/X sky130_fd_sc_hd__buf_1
X_4236_ _4236_/A VGND VGND VPWR VPWR _4236_/Y sky130_fd_sc_hd__inv_2
X_4167_ _3673_/B _5004_/Q _4166_/Y VGND VGND VPWR VPWR _4168_/A sky130_fd_sc_hd__o21ai_1
XFILLER_67_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3118_ _5081_/Q _3011_/X _3339_/A _3117_/Y VGND VGND VPWR VPWR _3119_/A sky130_fd_sc_hd__o22a_1
X_4098_ _4977_/Q VGND VGND VPWR VPWR _4099_/B sky130_fd_sc_hd__inv_2
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3049_ _5110_/Q VGND VGND VPWR VPWR _3049_/Y sky130_fd_sc_hd__inv_2
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2420_ _2426_/A _4659_/Y VGND VGND VPWR VPWR _2420_/X sky130_fd_sc_hd__or2_1
X_5070_ _3450_/X _5070_/D VGND VGND VPWR VPWR _5070_/Q sky130_fd_sc_hd__dfxtp_1
X_4021_ _3677_/B _5002_/Q _3677_/B _5002_/Q VGND VGND VPWR VPWR _4175_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4923_ _5028_/CLK _4923_/D VGND VGND VPWR VPWR _4923_/Q sky130_fd_sc_hd__dfxtp_1
X_4854_ _5047_/CLK _4854_/D VGND VGND VPWR VPWR _4854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4785_ _5139_/Q _4785_/D VGND VGND VPWR VPWR _4785_/Q sky130_fd_sc_hd__dfxtp_1
X_3805_ _3630_/B _5024_/Q _4913_/Q _3804_/Y VGND VGND VPWR VPWR _3806_/A sky130_fd_sc_hd__o22a_1
X_3736_ _3736_/A _3736_/B VGND VGND VPWR VPWR _4976_/D sky130_fd_sc_hd__nor2_1
X_3667_ _4895_/Q VGND VGND VPWR VPWR _3668_/B sky130_fd_sc_hd__inv_2
X_3598_ _4926_/Q VGND VGND VPWR VPWR _3599_/B sky130_fd_sc_hd__inv_2
X_2618_ _4948_/Q VGND VGND VPWR VPWR _2680_/A sky130_fd_sc_hd__clkbuf_2
X_2549_ _4722_/Y _2548_/Y _4728_/A VGND VGND VPWR VPWR _2549_/Y sky130_fd_sc_hd__o21ai_1
X_4219_ _4219_/A VGND VGND VPWR VPWR _4219_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4570_ _4569_/A _4568_/Y _4569_/Y _4568_/A _4539_/X VGND VGND VPWR VPWR _4874_/D
+ sky130_fd_sc_hd__o221a_1
X_3521_ input1/X input8/X VGND VGND VPWR VPWR _3522_/B sky130_fd_sc_hd__or2_1
X_3452_ _5070_/Q _3451_/Y _3435_/X _3452_/C1 VGND VGND VPWR VPWR _5070_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3383_ _3351_/A _3383_/A2 _3371_/X _3380_/Y VGND VGND VPWR VPWR _5093_/D sky130_fd_sc_hd__a211oi_1
X_2403_ _4657_/Y _4659_/Y _2426_/A _2402_/X VGND VGND VPWR VPWR _2416_/A sky130_fd_sc_hd__o31a_1
X_5122_ _3226_/X _5122_/D VGND VGND VPWR VPWR _5122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5053_ _5139_/CLK _5053_/D VGND VGND VPWR VPWR _5053_/Q sky130_fd_sc_hd__dfxtp_1
X_4004_ _4004_/A VGND VGND VPWR VPWR _4004_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4906_ _5018_/CLK _4906_/D VGND VGND VPWR VPWR _4906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4837_ _5028_/CLK _4837_/D VGND VGND VPWR VPWR _4837_/Q sky130_fd_sc_hd__dfxtp_1
X_4768_ _2820_/X _2811_/X _4770_/S VGND VGND VPWR VPWR _4785_/D sky130_fd_sc_hd__mux2_2
X_4699_ _4434_/A _3025_/A _4802_/Q _5115_/Q VGND VGND VPWR VPWR _4700_/B sky130_fd_sc_hd__o22a_1
X_3719_ _3725_/A _3719_/B VGND VGND VPWR VPWR _4984_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2952_ _5130_/Q VGND VGND VPWR VPWR _2952_/X sky130_fd_sc_hd__clkbuf_2
X_2883_ _2881_/Y _2882_/Y _3518_/B VGND VGND VPWR VPWR _2885_/A sky130_fd_sc_hd__o21ai_2
X_4622_ _4626_/A _4622_/B VGND VGND VPWR VPWR _4847_/D sky130_fd_sc_hd__nor2_1
X_4553_ _4630_/B _4840_/Q _4552_/Y VGND VGND VPWR VPWR _4554_/A sky130_fd_sc_hd__o21ai_1
X_4484_ _4484_/A VGND VGND VPWR VPWR _4484_/Y sky130_fd_sc_hd__inv_2
X_3504_ _3501_/Y _3502_/Y _3503_/X VGND VGND VPWR VPWR _3504_/X sky130_fd_sc_hd__o21a_1
X_3435_ _3978_/A VGND VGND VPWR VPWR _3435_/X sky130_fd_sc_hd__clkbuf_2
X_3366_ _3366_/A VGND VGND VPWR VPWR _3366_/Y sky130_fd_sc_hd__inv_2
X_5105_ _3305_/X _5105_/D VGND VGND VPWR VPWR _5105_/Q sky130_fd_sc_hd__dfxtp_1
X_3297_ _3312_/A VGND VGND VPWR VPWR _3297_/X sky130_fd_sc_hd__buf_1
X_5036_ _5047_/CLK _5036_/D VGND VGND VPWR VPWR _5036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput23 _4785_/Q VGND VGND VPWR VPWR DATA[13] sky130_fd_sc_hd__clkbuf_2
Xoutput34 _4781_/Q VGND VGND VPWR VPWR DATA[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3220_ _3220_/A VGND VGND VPWR VPWR _3220_/Y sky130_fd_sc_hd__inv_2
X_3151_ _3151_/A VGND VGND VPWR VPWR _3151_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3082_ _5067_/Q _5104_/Q _3081_/Y VGND VGND VPWR VPWR _3083_/A sky130_fd_sc_hd__a21oi_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3984_ _3984_/A _3984_/B VGND VGND VPWR VPWR _3985_/C sky130_fd_sc_hd__nand2_1
X_2935_ _5098_/Q VGND VGND VPWR VPWR _3356_/A sky130_fd_sc_hd__clkinvlp_4
X_2866_ _2866_/A _3503_/B VGND VGND VPWR VPWR _3512_/B sky130_fd_sc_hd__nor2_4
X_4605_ _4608_/A _4605_/B VGND VGND VPWR VPWR _4861_/D sky130_fd_sc_hd__nor2_1
X_2797_ _4968_/Q _2781_/X _2796_/X VGND VGND VPWR VPWR _2800_/C sky130_fd_sc_hd__o21a_1
X_4536_ _4536_/A _4536_/B VGND VGND VPWR VPWR _4536_/Y sky130_fd_sc_hd__nand2_1
X_4467_ _4821_/Q VGND VGND VPWR VPWR _4607_/B sky130_fd_sc_hd__inv_2
X_3418_ _5082_/Q _3417_/Y _3406_/X _3418_/C1 VGND VGND VPWR VPWR _5082_/D sky130_fd_sc_hd__o211a_1
X_4398_ _4722_/A _4830_/Q VGND VGND VPWR VPWR _4398_/Y sky130_fd_sc_hd__nor2_4
X_3349_ _3349_/A _3349_/B VGND VGND VPWR VPWR _3350_/B sky130_fd_sc_hd__or2_1
X_5019_ _5028_/CLK _5019_/D VGND VGND VPWR VPWR _5019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2720_ _2720_/A _2720_/B _2720_/C _2720_/D VGND VGND VPWR VPWR _2720_/X sky130_fd_sc_hd__or4_4
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2651_ _2791_/A VGND VGND VPWR VPWR _2651_/X sky130_fd_sc_hd__clkbuf_2
X_2582_ _2582_/A VGND VGND VPWR VPWR _2772_/A sky130_fd_sc_hd__inv_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4321_ _4849_/Q VGND VGND VPWR VPWR _4322_/B sky130_fd_sc_hd__inv_2
X_4252_ _4252_/A VGND VGND VPWR VPWR _4255_/A sky130_fd_sc_hd__inv_2
X_3203_ _3225_/A VGND VGND VPWR VPWR _3222_/A sky130_fd_sc_hd__buf_1
XFILLER_79_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4183_ _4183_/A VGND VGND VPWR VPWR _4183_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3134_ _5089_/Q _2977_/X _3133_/X VGND VGND VPWR VPWR _3134_/Y sky130_fd_sc_hd__o21ai_1
X_3065_ _3328_/A _3064_/X _5070_/Q _5107_/Q VGND VGND VPWR VPWR _3292_/A sky130_fd_sc_hd__o22a_1
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3967_ _3967_/A VGND VGND VPWR VPWR _3967_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2918_ _3485_/A _2879_/A _5059_/Q _2879_/Y _2917_/X VGND VGND VPWR VPWR _2918_/X
+ sky130_fd_sc_hd__o221a_1
X_3898_ _3766_/A _3905_/B _3868_/Y VGND VGND VPWR VPWR _3899_/B sky130_fd_sc_hd__o21ai_1
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2849_ _2881_/A _2882_/A VGND VGND VPWR VPWR _3518_/B sky130_fd_sc_hd__or2_2
X_4519_ _4546_/A _4450_/A _4351_/B VGND VGND VPWR VPWR _4520_/A sky130_fd_sc_hd__o21ai_1
XFILLER_58_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4870_ _5018_/CLK _4870_/D VGND VGND VPWR VPWR _4870_/Q sky130_fd_sc_hd__dfxtp_1
X_3821_ _4907_/Q _3820_/B _3820_/Y VGND VGND VPWR VPWR _3822_/A sky130_fd_sc_hd__a21oi_2
X_3752_ _4933_/Q _3751_/B _3751_/Y VGND VGND VPWR VPWR _3753_/A sky130_fd_sc_hd__a21oi_2
X_3683_ _3692_/A _3683_/B VGND VGND VPWR VPWR _5000_/D sky130_fd_sc_hd__nor2_1
X_2703_ _2703_/A _2756_/B VGND VGND VPWR VPWR _2703_/X sky130_fd_sc_hd__or2_1
X_2634_ _2666_/A _4958_/Q VGND VGND VPWR VPWR _2637_/B sky130_fd_sc_hd__or2b_1
X_2565_ _4945_/Q VGND VGND VPWR VPWR _2636_/B sky130_fd_sc_hd__clkbuf_2
X_4304_ _4488_/A _4304_/B VGND VGND VPWR VPWR _4305_/B sky130_fd_sc_hd__or2_1
X_2496_ _4752_/Y _2494_/Y _4752_/A _2494_/A _2495_/X VGND VGND VPWR VPWR _4805_/D
+ sky130_fd_sc_hd__o221a_1
X_4235_ _4074_/A _4234_/Y _4072_/A _4234_/A _4229_/X VGND VGND VPWR VPWR _4913_/D
+ sky130_fd_sc_hd__o221a_1
X_4166_ _4166_/A _4166_/B VGND VGND VPWR VPWR _4166_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3117_ _5118_/Q VGND VGND VPWR VPWR _3117_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4097_ _4097_/A _4260_/B VGND VGND VPWR VPWR _4111_/C sky130_fd_sc_hd__nand2_1
XFILLER_55_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3048_ _5073_/Q VGND VGND VPWR VPWR _3331_/A sky130_fd_sc_hd__clkinv_1
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4999_ _5047_/CLK _4999_/D VGND VGND VPWR VPWR _4999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4020_ _3668_/B _5006_/Q _3668_/B _5006_/Q VGND VGND VPWR VPWR _4160_/B sky130_fd_sc_hd__a2bb2o_1
X_4922_ _5028_/CLK _4922_/D VGND VGND VPWR VPWR _4922_/Q sky130_fd_sc_hd__dfxtp_1
X_4853_ _5047_/CLK _4853_/D VGND VGND VPWR VPWR _4853_/Q sky130_fd_sc_hd__dfxtp_1
X_4784_ _5047_/CLK _4784_/D VGND VGND VPWR VPWR _4784_/Q sky130_fd_sc_hd__dfxtp_1
X_3804_ _5024_/Q VGND VGND VPWR VPWR _3804_/Y sky130_fd_sc_hd__inv_2
X_3735_ _4865_/Q VGND VGND VPWR VPWR _3736_/B sky130_fd_sc_hd__inv_2
X_3666_ _3668_/A _3666_/B VGND VGND VPWR VPWR _5007_/D sky130_fd_sc_hd__nor2_1
X_3597_ _3599_/A _3597_/B VGND VGND VPWR VPWR _5038_/D sky130_fd_sc_hd__nor2_1
X_2617_ _2721_/A _2787_/A VGND VGND VPWR VPWR _2617_/Y sky130_fd_sc_hd__nor2_1
X_2548_ _2548_/A VGND VGND VPWR VPWR _2548_/Y sky130_fd_sc_hd__inv_2
X_2479_ _3459_/A VGND VGND VPWR VPWR _2497_/A sky130_fd_sc_hd__buf_1
X_4218_ _4126_/A _4217_/Y _4123_/A _4217_/A _4190_/X VGND VGND VPWR VPWR _4917_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4149_ _3664_/B _5008_/Q _4155_/B VGND VGND VPWR VPWR _4150_/A sky130_fd_sc_hd__o21ai_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3520_ _5055_/Q _3519_/X _5055_/Q _3519_/X VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3451_ _3451_/A VGND VGND VPWR VPWR _3451_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3382_ _3382_/A VGND VGND VPWR VPWR _3382_/X sky130_fd_sc_hd__buf_1
X_2402_ _4608_/B _2945_/X _4655_/Y _4607_/B _3143_/Y VGND VGND VPWR VPWR _2402_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5121_ _3231_/X _5121_/D VGND VGND VPWR VPWR _5121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5052_ _5139_/CLK _5052_/D VGND VGND VPWR VPWR _5052_/Q sky130_fd_sc_hd__dfxtp_1
X_4003_ _3835_/Y _4002_/Y _3835_/A _4002_/A _3976_/X VGND VGND VPWR VPWR _4940_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_65_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4905_ _5018_/CLK _4905_/D VGND VGND VPWR VPWR _4905_/Q sky130_fd_sc_hd__dfxtp_1
X_4836_ _5028_/CLK _4836_/D VGND VGND VPWR VPWR _4836_/Q sky130_fd_sc_hd__dfxtp_1
X_4767_ _2810_/X _2801_/X _4770_/S VGND VGND VPWR VPWR _4784_/D sky130_fd_sc_hd__mux2_2
X_4698_ _4803_/Q _5116_/Q _4697_/Y VGND VGND VPWR VPWR _4700_/A sky130_fd_sc_hd__a21oi_2
X_3718_ _4873_/Q VGND VGND VPWR VPWR _3719_/B sky130_fd_sc_hd__inv_2
X_3649_ _4904_/Q VGND VGND VPWR VPWR _3825_/A sky130_fd_sc_hd__inv_2
XFILLER_75_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2951_ _2951_/A VGND VGND VPWR VPWR _3189_/A sky130_fd_sc_hd__inv_2
X_2882_ _2882_/A VGND VGND VPWR VPWR _2882_/Y sky130_fd_sc_hd__inv_2
X_4621_ _4621_/A VGND VGND VPWR VPWR _4626_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4552_ _4552_/A _4552_/B VGND VGND VPWR VPWR _4552_/Y sky130_fd_sc_hd__nand2_1
X_4483_ _4608_/B _4858_/Q _4487_/B VGND VGND VPWR VPWR _4484_/A sky130_fd_sc_hd__o21ai_1
X_3503_ _3508_/A _3503_/B VGND VGND VPWR VPWR _3503_/X sky130_fd_sc_hd__or2_1
X_3434_ _3434_/A VGND VGND VPWR VPWR _3434_/Y sky130_fd_sc_hd__inv_2
X_3365_ _3365_/A VGND VGND VPWR VPWR _3365_/X sky130_fd_sc_hd__buf_1
X_3296_ _3368_/A VGND VGND VPWR VPWR _3312_/A sky130_fd_sc_hd__buf_1
X_5104_ _3307_/X _5104_/D VGND VGND VPWR VPWR _5104_/Q sky130_fd_sc_hd__dfxtp_2
X_5035_ _5047_/CLK _5035_/D VGND VGND VPWR VPWR _5035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4819_ _2428_/X _4819_/D VGND VGND VPWR VPWR _4819_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput24 _4786_/Q VGND VGND VPWR VPWR DATA[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput35 _4825_/Q VGND VGND VPWR VPWR data_en sky130_fd_sc_hd__clkbuf_2
XFILLER_29_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3150_ _3150_/A VGND VGND VPWR VPWR _3150_/Y sky130_fd_sc_hd__inv_2
X_3081_ _5067_/Q _5104_/Q VGND VGND VPWR VPWR _3081_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3983_ _3817_/A _3982_/Y _3815_/A _3982_/A _3976_/X VGND VGND VPWR VPWR _4946_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2934_ _2934_/A VGND VGND VPWR VPWR _2934_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2865_ input2/X VGND VGND VPWR VPWR _2866_/A sky130_fd_sc_hd__buf_2
X_4604_ _4608_/A _4604_/B VGND VGND VPWR VPWR _4862_/D sky130_fd_sc_hd__nor2_1
X_2796_ _2796_/A VGND VGND VPWR VPWR _2796_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4535_ _4546_/A _4446_/B _4347_/Y VGND VGND VPWR VPWR _4536_/B sky130_fd_sc_hd__o21ai_1
X_4466_ _4466_/A VGND VGND VPWR VPWR _4608_/B sky130_fd_sc_hd__clkbuf_2
X_3417_ _3417_/A VGND VGND VPWR VPWR _3417_/Y sky130_fd_sc_hd__clkinvlp_2
X_4397_ _4792_/Q VGND VGND VPWR VPWR _4722_/A sky130_fd_sc_hd__clkinv_4
X_3348_ _3348_/A _3348_/B VGND VGND VPWR VPWR _3349_/B sky130_fd_sc_hd__or2_1
X_3279_ _3274_/A _3274_/B _3258_/X _3274_/Y VGND VGND VPWR VPWR _5111_/D sky130_fd_sc_hd__o211a_1
XFILLER_26_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5018_ _5018_/CLK _5018_/D VGND VGND VPWR VPWR _5018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2650_ _2650_/A VGND VGND VPWR VPWR _2791_/A sky130_fd_sc_hd__inv_2
X_2581_ _2911_/Y _3517_/A _3516_/B _2584_/B VGND VGND VPWR VPWR _2582_/A sky130_fd_sc_hd__or4_4
X_4320_ _4320_/A _4320_/B VGND VGND VPWR VPWR _4320_/X sky130_fd_sc_hd__or2_1
X_4251_ _4481_/A _4251_/B _4251_/C VGND VGND VPWR VPWR _4908_/D sky130_fd_sc_hd__and3_1
X_3202_ _3201_/A _3201_/B _3186_/X _3201_/Y VGND VGND VPWR VPWR _5128_/D sky130_fd_sc_hd__o211a_1
X_4182_ _3683_/B _5000_/Q _4181_/Y VGND VGND VPWR VPWR _4183_/A sky130_fd_sc_hd__o21ai_1
X_3133_ _5089_/Q _2977_/X _5088_/Q _5125_/Q VGND VGND VPWR VPWR _3133_/X sky130_fd_sc_hd__a22o_1
X_3064_ _3064_/A VGND VGND VPWR VPWR _3064_/X sky130_fd_sc_hd__clkbuf_2
X_3966_ _3808_/A _3965_/Y _3806_/A _3965_/A _3936_/X VGND VGND VPWR VPWR _4950_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2917_ _3481_/A _2872_/Y _2887_/X _2916_/X VGND VGND VPWR VPWR _2917_/X sky130_fd_sc_hd__o211a_1
XFILLER_31_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3897_ _3897_/A VGND VGND VPWR VPWR _3905_/B sky130_fd_sc_hd__inv_2
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2848_ _2891_/A _2848_/B VGND VGND VPWR VPWR _2882_/A sky130_fd_sc_hd__or2_1
X_2779_ _2811_/A _2777_/X _2778_/X VGND VGND VPWR VPWR _2780_/D sky130_fd_sc_hd__o21a_1
X_4518_ _4578_/A _4518_/B _4518_/C VGND VGND VPWR VPWR _4887_/D sky130_fd_sc_hd__and3_1
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4449_ _4326_/A _4848_/Q _4325_/A _4848_/Q VGND VGND VPWR VPWR _4522_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3820_ _4907_/Q _3820_/B VGND VGND VPWR VPWR _3820_/Y sky130_fd_sc_hd__nor2_1
X_3751_ _4933_/Q _3751_/B VGND VGND VPWR VPWR _3751_/Y sky130_fd_sc_hd__nor2_1
X_2702_ _2831_/B VGND VGND VPWR VPWR _2756_/B sky130_fd_sc_hd__buf_1
XFILLER_9_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3682_ _4889_/Q VGND VGND VPWR VPWR _3683_/B sky130_fd_sc_hd__inv_2
X_2633_ _4947_/Q VGND VGND VPWR VPWR _2666_/A sky130_fd_sc_hd__clkbuf_2
X_2564_ _4735_/A _3096_/B _4788_/Q _5101_/Q _3985_/A VGND VGND VPWR VPWR _4788_/D
+ sky130_fd_sc_hd__o221a_1
X_4303_ _4303_/A VGND VGND VPWR VPWR _4304_/B sky130_fd_sc_hd__inv_2
X_2495_ _4575_/A VGND VGND VPWR VPWR _2495_/X sky130_fd_sc_hd__buf_2
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4234_ _4234_/A VGND VGND VPWR VPWR _4234_/Y sky130_fd_sc_hd__inv_2
X_4165_ _4032_/A _4171_/B _4134_/Y VGND VGND VPWR VPWR _4166_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3116_ _5081_/Q VGND VGND VPWR VPWR _3339_/A sky130_fd_sc_hd__inv_2
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ _4091_/A _4978_/Q _4091_/Y VGND VGND VPWR VPWR _4260_/B sky130_fd_sc_hd__a21oi_4
X_3047_ _3276_/A _3274_/A VGND VGND VPWR VPWR _3058_/A sky130_fd_sc_hd__nand2_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4998_ _5047_/CLK _4998_/D VGND VGND VPWR VPWR _4998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3949_ _3622_/B _5027_/Q _3948_/X VGND VGND VPWR VPWR _3950_/A sky130_fd_sc_hd__o21ai_1
XFILLER_48_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4921_ _5047_/CLK _4921_/D VGND VGND VPWR VPWR _4921_/Q sky130_fd_sc_hd__dfxtp_1
X_4852_ _5047_/CLK _4852_/D VGND VGND VPWR VPWR _4852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3803_ _3803_/A _3954_/A VGND VGND VPWR VPWR _3809_/A sky130_fd_sc_hd__or2_1
X_4783_ _5018_/CLK _4783_/D VGND VGND VPWR VPWR _4783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3734_ _3736_/A _3734_/B VGND VGND VPWR VPWR _4977_/D sky130_fd_sc_hd__nor2_1
X_3665_ _4896_/Q VGND VGND VPWR VPWR _3666_/B sky130_fd_sc_hd__inv_2
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2616_ _2616_/A _2616_/B _2616_/C VGND VGND VPWR VPWR _2787_/A sky130_fd_sc_hd__nor3_4
X_3596_ _4927_/Q VGND VGND VPWR VPWR _3597_/B sky130_fd_sc_hd__inv_2
X_2547_ _2547_/A _4728_/B VGND VGND VPWR VPWR _2548_/A sky130_fd_sc_hd__nand2_1
X_2478_ _4684_/A _2477_/Y _4681_/A _2477_/A _2423_/X VGND VGND VPWR VPWR _4809_/D
+ sky130_fd_sc_hd__o221a_1
X_4217_ _4217_/A VGND VGND VPWR VPWR _4217_/Y sky130_fd_sc_hd__inv_2
X_4148_ _4154_/A _4154_/B VGND VGND VPWR VPWR _4155_/B sky130_fd_sc_hd__or2_1
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4079_ _4983_/Q VGND VGND VPWR VPWR _4079_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3450_ _3455_/A VGND VGND VPWR VPWR _3450_/X sky130_fd_sc_hd__buf_1
X_3381_ _5094_/Q _3380_/Y _3375_/X _3381_/C1 VGND VGND VPWR VPWR _5094_/D sky130_fd_sc_hd__o211a_1
X_2401_ _4669_/X _4678_/X _2462_/A _2400_/X VGND VGND VPWR VPWR _2426_/A sky130_fd_sc_hd__o31a_1
X_5120_ _3233_/X _5120_/D VGND VGND VPWR VPWR _5120_/Q sky130_fd_sc_hd__dfxtp_1
X_5051_ _5063_/CLK _5051_/D VGND VGND VPWR VPWR _5051_/Q sky130_fd_sc_hd__dfxtp_1
X_4002_ _4002_/A VGND VGND VPWR VPWR _4002_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4904_ _5018_/CLK _4904_/D VGND VGND VPWR VPWR _4904_/Q sky130_fd_sc_hd__dfxtp_1
X_4835_ _5028_/CLK _4835_/D VGND VGND VPWR VPWR _4835_/Q sky130_fd_sc_hd__dfxtp_1
X_4766_ _2800_/X _2786_/X _4770_/S VGND VGND VPWR VPWR _4783_/D sky130_fd_sc_hd__mux2_1
X_3717_ _3725_/A _3717_/B VGND VGND VPWR VPWR _4985_/D sky130_fd_sc_hd__nor2_1
X_4697_ _4803_/Q _5116_/Q VGND VGND VPWR VPWR _4697_/Y sky130_fd_sc_hd__nor2_1
X_3648_ _3656_/A _3824_/A VGND VGND VPWR VPWR _5016_/D sky130_fd_sc_hd__nor2_1
X_3579_ _4935_/Q VGND VGND VPWR VPWR _3580_/B sky130_fd_sc_hd__inv_2
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2950_ _5092_/Q _5129_/Q _3350_/A _2949_/Y VGND VGND VPWR VPWR _2951_/A sky130_fd_sc_hd__o22a_1
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2881_ _2881_/A VGND VGND VPWR VPWR _2881_/Y sky130_fd_sc_hd__inv_2
X_4620_ _4620_/A _4620_/B VGND VGND VPWR VPWR _4848_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4551_ _4372_/B _4557_/B _4427_/Y VGND VGND VPWR VPWR _4552_/B sky130_fd_sc_hd__o21ai_1
X_4482_ _4486_/A _4486_/B VGND VGND VPWR VPWR _4487_/B sky130_fd_sc_hd__or2_1
X_3502_ _3508_/A _3502_/B VGND VGND VPWR VPWR _3502_/Y sky130_fd_sc_hd__nor2_1
X_3433_ _3442_/A VGND VGND VPWR VPWR _3433_/X sky130_fd_sc_hd__buf_1
X_5103_ _3312_/X _5103_/D VGND VGND VPWR VPWR _5103_/Q sky130_fd_sc_hd__dfxtp_1
X_3364_ _3357_/A _3364_/A2 _4647_/A _3358_/Y VGND VGND VPWR VPWR _5099_/D sky130_fd_sc_hd__a211oi_2
X_3295_ _3103_/A _3294_/Y _3061_/A _3294_/A _3267_/X VGND VGND VPWR VPWR _5108_/D
+ sky130_fd_sc_hd__o221a_1
X_5034_ _5047_/CLK _5034_/D VGND VGND VPWR VPWR _5034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4818_ _2437_/X _4818_/D VGND VGND VPWR VPWR _4818_/Q sky130_fd_sc_hd__dfxtp_1
X_4749_ _4706_/A _4743_/Y _4706_/X _4747_/X _4748_/X VGND VGND VPWR VPWR _4749_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput25 _4787_/Q VGND VGND VPWR VPWR DATA[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_29_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3080_ _3080_/A _3300_/B VGND VGND VPWR VPWR _3103_/C sky130_fd_sc_hd__nand2_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3982_ _3982_/A VGND VGND VPWR VPWR _3982_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2933_ _5099_/Q _5136_/Q _2932_/Y VGND VGND VPWR VPWR _2934_/A sky130_fd_sc_hd__a21oi_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2864_ input3/X VGND VGND VPWR VPWR _2864_/Y sky130_fd_sc_hd__inv_2
X_2795_ _2795_/A _2795_/B _2795_/C _2795_/D VGND VGND VPWR VPWR _2800_/B sky130_fd_sc_hd__or4_4
X_4603_ _4824_/Q VGND VGND VPWR VPWR _4604_/B sky130_fd_sc_hd__inv_2
X_4534_ _4534_/A VGND VGND VPWR VPWR _4536_/A sky130_fd_sc_hd__inv_2
X_4465_ _4305_/X _4320_/X _4517_/A _4464_/X VGND VGND VPWR VPWR _4486_/A sky130_fd_sc_hd__o31a_1
X_3416_ _3426_/A VGND VGND VPWR VPWR _3416_/X sky130_fd_sc_hd__buf_1
X_4396_ _4396_/A _4831_/Q VGND VGND VPWR VPWR _4396_/Y sky130_fd_sc_hd__nor2_2
X_3347_ _3347_/A _3347_/B VGND VGND VPWR VPWR _3348_/B sky130_fd_sc_hd__or2_1
X_3278_ _3289_/A VGND VGND VPWR VPWR _3278_/X sky130_fd_sc_hd__buf_1
X_5017_ _5018_/CLK _5017_/D VGND VGND VPWR VPWR _5017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2580_ _2881_/A _2580_/B VGND VGND VPWR VPWR _2584_/B sky130_fd_sc_hd__or2_1
X_4250_ _4250_/A _4250_/B VGND VGND VPWR VPWR _4251_/C sky130_fd_sc_hd__nand2_1
XFILLER_79_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4181_ _4181_/A _4181_/B VGND VGND VPWR VPWR _4181_/Y sky130_fd_sc_hd__nand2_1
X_3201_ _3201_/A _3201_/B VGND VGND VPWR VPWR _3201_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3132_ _5093_/Q _2952_/X _3131_/X VGND VGND VPWR VPWR _3132_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3063_ _5107_/Q VGND VGND VPWR VPWR _3064_/A sky130_fd_sc_hd__inv_2
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3965_ _3965_/A VGND VGND VPWR VPWR _3965_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3896_ _3923_/A _3775_/X _3872_/X VGND VGND VPWR VPWR _3897_/A sky130_fd_sc_hd__o21ai_2
X_2916_ _5055_/Q _2889_/Y _3480_/A _2889_/A _2915_/Y VGND VGND VPWR VPWR _2916_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2847_ _3516_/A _3515_/B VGND VGND VPWR VPWR _2848_/B sky130_fd_sc_hd__or2_2
X_2778_ _2778_/A VGND VGND VPWR VPWR _2778_/X sky130_fd_sc_hd__buf_1
X_4517_ _4517_/A _4517_/B VGND VGND VPWR VPWR _4518_/C sky130_fd_sc_hd__nand2_1
X_4448_ _4448_/A VGND VGND VPWR VPWR _4450_/B sky130_fd_sc_hd__inv_2
X_4379_ _4797_/Q VGND VGND VPWR VPWR _4379_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ _5044_/Q VGND VGND VPWR VPWR _3751_/B sky130_fd_sc_hd__inv_2
XFILLER_20_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2701_ _2701_/A _2701_/B _2701_/C _2701_/D VGND VGND VPWR VPWR _2701_/X sky130_fd_sc_hd__or4_1
X_3681_ _3726_/A VGND VGND VPWR VPWR _3692_/A sky130_fd_sc_hd__clkbuf_2
X_2632_ _4951_/Q _2632_/B _2632_/C _2632_/D VGND VGND VPWR VPWR _2650_/A sky130_fd_sc_hd__or4_4
X_2563_ _3225_/A VGND VGND VPWR VPWR _2563_/X sky130_fd_sc_hd__buf_1
X_4302_ _4819_/Q _4301_/B _4301_/Y VGND VGND VPWR VPWR _4303_/A sky130_fd_sc_hd__a21oi_2
X_2494_ _2494_/A VGND VGND VPWR VPWR _2494_/Y sky130_fd_sc_hd__inv_2
X_4233_ _3714_/B _4986_/Q _4232_/X VGND VGND VPWR VPWR _4234_/A sky130_fd_sc_hd__o21ai_1
X_4164_ _4164_/A VGND VGND VPWR VPWR _4171_/B sky130_fd_sc_hd__inv_2
X_3115_ _3038_/X _3058_/X _3286_/A _3114_/X VGND VGND VPWR VPWR _3250_/A sky130_fd_sc_hd__o31a_2
X_4095_ _4090_/A _4979_/Q _4090_/Y VGND VGND VPWR VPWR _4097_/A sky130_fd_sc_hd__a21oi_2
X_3046_ _3332_/A _3045_/X _5074_/Q _5111_/Q VGND VGND VPWR VPWR _3274_/A sky130_fd_sc_hd__o22a_1
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4997_ _5028_/CLK _4997_/D VGND VGND VPWR VPWR _4997_/Q sky130_fd_sc_hd__dfxtp_1
X_3948_ _3952_/A _3948_/B VGND VGND VPWR VPWR _3948_/X sky130_fd_sc_hd__or2_1
X_3879_ _3748_/Y _3887_/B _3887_/A _3878_/X VGND VGND VPWR VPWR _3880_/A sky130_fd_sc_hd__o31a_1
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4920_ _5047_/CLK _4920_/D VGND VGND VPWR VPWR _4920_/Q sky130_fd_sc_hd__dfxtp_1
X_4851_ _5047_/CLK _4851_/D VGND VGND VPWR VPWR _4851_/Q sky130_fd_sc_hd__dfxtp_1
X_3802_ _3628_/B _5025_/Q _3628_/B _5025_/Q VGND VGND VPWR VPWR _3954_/A sky130_fd_sc_hd__a2bb2o_1
X_4782_ _5018_/CLK _4782_/D VGND VGND VPWR VPWR _4782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3733_ _4866_/Q VGND VGND VPWR VPWR _3734_/B sky130_fd_sc_hd__inv_2
X_3664_ _3668_/A _3664_/B VGND VGND VPWR VPWR _5008_/D sky130_fd_sc_hd__nor2_1
X_2615_ _4956_/Q _4955_/Q _2615_/C _4967_/Q VGND VGND VPWR VPWR _2616_/B sky130_fd_sc_hd__or4b_4
X_3595_ _3599_/A _3595_/B VGND VGND VPWR VPWR _5039_/D sky130_fd_sc_hd__nor2_1
X_2546_ _2560_/A VGND VGND VPWR VPWR _2546_/X sky130_fd_sc_hd__buf_1
X_2477_ _2477_/A VGND VGND VPWR VPWR _2477_/Y sky130_fd_sc_hd__inv_2
X_4216_ _3706_/B _4990_/Q _4215_/X VGND VGND VPWR VPWR _4217_/A sky130_fd_sc_hd__o21ai_1
X_4147_ _4010_/Y _4146_/A _4010_/A _4146_/Y _3976_/X VGND VGND VPWR VPWR _4936_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4078_ _4243_/A _4238_/A VGND VGND VPWR VPWR _4084_/A sky130_fd_sc_hd__or2_1
XFILLER_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3029_ _5114_/Q VGND VGND VPWR VPWR _3029_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2400_ _4669_/B _2394_/Y _4669_/X _2398_/X _2399_/X VGND VGND VPWR VPWR _2400_/X
+ sky130_fd_sc_hd__o221a_1
X_3380_ _3380_/A VGND VGND VPWR VPWR _3380_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5050_ _5063_/CLK _5050_/D VGND VGND VPWR VPWR _5050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4001_ _3654_/B _5013_/Q _4000_/X VGND VGND VPWR VPWR _4002_/A sky130_fd_sc_hd__o21ai_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4903_ _5018_/CLK _4903_/D VGND VGND VPWR VPWR _4903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4834_ _5028_/CLK _4834_/D VGND VGND VPWR VPWR _4834_/Q sky130_fd_sc_hd__dfxtp_1
X_4765_ _2785_/X _2768_/X _4770_/S VGND VGND VPWR VPWR _4782_/D sky130_fd_sc_hd__mux2_1
X_3716_ _4874_/Q VGND VGND VPWR VPWR _3717_/B sky130_fd_sc_hd__inv_2
X_4696_ _4619_/B _2988_/Y _4620_/B _2991_/X _4695_/X VGND VGND VPWR VPWR _4696_/X
+ sky130_fd_sc_hd__o221a_1
X_3647_ _4905_/Q VGND VGND VPWR VPWR _3824_/A sky130_fd_sc_hd__inv_2
X_3578_ _3612_/A VGND VGND VPWR VPWR _3588_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2529_ _4741_/X _4714_/B VGND VGND VPWR VPWR _2529_/X sky130_fd_sc_hd__or2_1
XFILLER_29_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2880_ _5063_/Q VGND VGND VPWR VPWR _2880_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4550_ _4550_/A VGND VGND VPWR VPWR _4557_/B sky130_fd_sc_hd__inv_2
X_4481_ _4481_/A _4481_/B _4481_/C VGND VGND VPWR VPWR _4897_/D sky130_fd_sc_hd__and3_1
X_3501_ _3501_/A VGND VGND VPWR VPWR _3501_/Y sky130_fd_sc_hd__inv_2
X_3432_ _3335_/A _3432_/A2 _3431_/X _3427_/Y VGND VGND VPWR VPWR _5077_/D sky130_fd_sc_hd__a211oi_1
X_3363_ _3737_/A VGND VGND VPWR VPWR _4647_/A sky130_fd_sc_hd__clkbuf_4
X_5102_ _3315_/X _5102_/D VGND VGND VPWR VPWR _5102_/Q sky130_fd_sc_hd__dfxtp_1
X_3294_ _3294_/A VGND VGND VPWR VPWR _3294_/Y sky130_fd_sc_hd__inv_2
X_5033_ _5047_/CLK _5033_/D VGND VGND VPWR VPWR _5033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4817_ _2439_/X _4817_/D VGND VGND VPWR VPWR _4817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4748_ _4630_/B _3025_/X _4697_/Y _4629_/B _3112_/Y VGND VGND VPWR VPWR _4748_/X
+ sky130_fd_sc_hd__o32a_1
X_4679_ _4811_/Q _5124_/Q VGND VGND VPWR VPWR _4679_/Y sky130_fd_sc_hd__nor2_2
Xoutput26 _4773_/Q VGND VGND VPWR VPWR DATA[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3981_ _3641_/B _5019_/Q _3985_/B VGND VGND VPWR VPWR _3982_/A sky130_fd_sc_hd__o21ai_1
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2932_ _5099_/Q _5136_/Q VGND VGND VPWR VPWR _2932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2863_ input5/X _3508_/B _3498_/B VGND VGND VPWR VPWR _2863_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2794_ _2821_/A _2777_/X _2778_/X VGND VGND VPWR VPWR _2795_/D sky130_fd_sc_hd__o21a_1
X_4602_ _4621_/A VGND VGND VPWR VPWR _4608_/A sky130_fd_sc_hd__clkbuf_2
X_4533_ _4532_/Y _4520_/A _4526_/X _4528_/X VGND VGND VPWR VPWR _4883_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4464_ _4305_/B _4454_/Y _4305_/X _4460_/X _4463_/X VGND VGND VPWR VPWR _4464_/X
+ sky130_fd_sc_hd__o221a_1
X_3415_ _3444_/A VGND VGND VPWR VPWR _3426_/A sky130_fd_sc_hd__buf_1
X_4395_ _4396_/A VGND VGND VPWR VPWR _4721_/A sky130_fd_sc_hd__buf_2
X_3346_ _3346_/A _3346_/B VGND VGND VPWR VPWR _3347_/B sky130_fd_sc_hd__or2_1
X_3277_ _3276_/A _3276_/B _3258_/X _3276_/Y VGND VGND VPWR VPWR _5112_/D sky130_fd_sc_hd__o211a_1
X_5016_ _5018_/CLK _5016_/D VGND VGND VPWR VPWR _5016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4180_ _4192_/A _4041_/B _4136_/Y VGND VGND VPWR VPWR _4181_/B sky130_fd_sc_hd__o21ai_1
X_3200_ _3348_/A _2972_/X _3199_/Y VGND VGND VPWR VPWR _3201_/B sky130_fd_sc_hd__o21ai_1
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3131_ _5092_/Q _5129_/Q _5093_/Q _2952_/X VGND VGND VPWR VPWR _3131_/X sky130_fd_sc_hd__a22o_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3062_ _5070_/Q VGND VGND VPWR VPWR _3328_/A sky130_fd_sc_hd__clkinvlp_4
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3964_ _3632_/B _5023_/Q _3963_/X VGND VGND VPWR VPWR _3965_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3895_ _3895_/A VGND VGND VPWR VPWR _3899_/A sky130_fd_sc_hd__inv_2
X_2915_ _5053_/Q _2894_/A _3478_/A _2894_/Y _2914_/X VGND VGND VPWR VPWR _2915_/Y
+ sky130_fd_sc_hd__a221oi_2
X_2846_ _3532_/A _2846_/B VGND VGND VPWR VPWR _3515_/B sky130_fd_sc_hd__or2_1
X_2777_ _2777_/A VGND VGND VPWR VPWR _2777_/X sky130_fd_sc_hd__buf_1
X_4516_ _4319_/A _4515_/Y _4315_/A _4515_/A _4501_/X VGND VGND VPWR VPWR _4888_/D
+ sky130_fd_sc_hd__o221a_1
X_4447_ _4811_/Q _4322_/B _4322_/Y VGND VGND VPWR VPWR _4448_/A sky130_fd_sc_hd__a21oi_2
X_4378_ _4797_/Q VGND VGND VPWR VPWR _4636_/B sky130_fd_sc_hd__inv_2
X_3329_ _3329_/A _3329_/B VGND VGND VPWR VPWR _3330_/B sky130_fd_sc_hd__or2_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2700_ _2811_/A _2613_/B _2663_/X VGND VGND VPWR VPWR _2701_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3680_ _3737_/A VGND VGND VPWR VPWR _3726_/A sky130_fd_sc_hd__buf_2
X_2631_ _2631_/A _4938_/Q _4937_/Q _4952_/Q VGND VGND VPWR VPWR _2632_/C sky130_fd_sc_hd__or4b_4
X_2562_ _2561_/X _4735_/X _3318_/C VGND VGND VPWR VPWR _4789_/D sky130_fd_sc_hd__and3b_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4301_ _4819_/Q _4301_/B VGND VGND VPWR VPWR _4301_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2493_ _4628_/B _3121_/Y _2492_/X VGND VGND VPWR VPWR _2494_/A sky130_fd_sc_hd__o21ai_1
X_4232_ _4236_/A _4232_/B VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__or2_1
X_4163_ _4192_/A _4041_/X _4138_/X VGND VGND VPWR VPWR _4164_/A sky130_fd_sc_hd__o21ai_1
X_3114_ _3038_/A _3106_/Y _3038_/X _3110_/X _3113_/X VGND VGND VPWR VPWR _3114_/X
+ sky130_fd_sc_hd__o221a_1
X_4094_ _3728_/B _4980_/Q _4086_/Y _3725_/B _4981_/Q VGND VGND VPWR VPWR _4094_/X
+ sky130_fd_sc_hd__o32a_1
X_3045_ _3045_/A VGND VGND VPWR VPWR _3045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4996_ _5028_/CLK _4996_/D VGND VGND VPWR VPWR _4996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3947_ _3943_/A _3943_/B _3939_/X _3943_/Y VGND VGND VPWR VPWR _4955_/D sky130_fd_sc_hd__o211a_1
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3878_ _3582_/B _5045_/Q _3746_/Y _3580_/B _5046_/Q VGND VGND VPWR VPWR _3878_/X
+ sky130_fd_sc_hd__o32a_1
X_2829_ _4968_/Q _2783_/X _2798_/X VGND VGND VPWR VPWR _2830_/D sky130_fd_sc_hd__o21a_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4850_ _5047_/CLK _4850_/D VGND VGND VPWR VPWR _4850_/Q sky130_fd_sc_hd__dfxtp_1
X_3801_ _3801_/A VGND VGND VPWR VPWR _3803_/A sky130_fd_sc_hd__inv_2
X_4781_ _5018_/CLK _4781_/D VGND VGND VPWR VPWR _4781_/Q sky130_fd_sc_hd__dfxtp_1
X_3732_ _3736_/A _4091_/A VGND VGND VPWR VPWR _4978_/D sky130_fd_sc_hd__nor2_1
X_3663_ _4897_/Q VGND VGND VPWR VPWR _3664_/B sky130_fd_sc_hd__inv_2
X_2614_ _4951_/Q VGND VGND VPWR VPWR _2721_/A sky130_fd_sc_hd__clkbuf_2
X_3594_ _4928_/Q VGND VGND VPWR VPWR _3595_/B sky130_fd_sc_hd__inv_2
X_2545_ _3384_/A VGND VGND VPWR VPWR _2560_/A sky130_fd_sc_hd__buf_1
X_2476_ _4623_/B _2998_/Y _2475_/X VGND VGND VPWR VPWR _2477_/A sky130_fd_sc_hd__o21ai_1
X_4215_ _4219_/A _4215_/B VGND VGND VPWR VPWR _4215_/X sky130_fd_sc_hd__or2_1
X_4146_ _4146_/A VGND VGND VPWR VPWR _4146_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ _3719_/B _4984_/Q _3719_/B _4984_/Q VGND VGND VPWR VPWR _4238_/A sky130_fd_sc_hd__a2bb2o_1
X_3028_ _5077_/Q VGND VGND VPWR VPWR _3335_/A sky130_fd_sc_hd__clkinv_1
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4979_ _5018_/CLK _4979_/D VGND VGND VPWR VPWR _4979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4000_ _4000_/A _4004_/A VGND VGND VPWR VPWR _4000_/X sky130_fd_sc_hd__or2_1
XFILLER_65_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _5018_/CLK _4902_/D VGND VGND VPWR VPWR _4902_/Q sky130_fd_sc_hd__dfxtp_1
X_4833_ _5139_/Q _4833_/D VGND VGND VPWR VPWR _4833_/Q sky130_fd_sc_hd__dfxtp_1
X_4764_ _2766_/X _2756_/X _4770_/S VGND VGND VPWR VPWR _4781_/D sky130_fd_sc_hd__mux2_1
X_3715_ _3726_/A VGND VGND VPWR VPWR _3725_/A sky130_fd_sc_hd__clkbuf_2
X_4695_ _4326_/A _2991_/A _4692_/X _4694_/Y VGND VGND VPWR VPWR _4695_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3646_ _3669_/A VGND VGND VPWR VPWR _3656_/A sky130_fd_sc_hd__clkbuf_2
X_3577_ _3660_/A _4936_/Q VGND VGND VPWR VPWR _5047_/D sky130_fd_sc_hd__and2_1
XFILLER_0_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2528_ _2543_/A VGND VGND VPWR VPWR _2528_/X sky130_fd_sc_hd__buf_1
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2459_ _2459_/A VGND VGND VPWR VPWR _2459_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4129_ _4129_/A VGND VGND VPWR VPWR _4131_/B sky130_fd_sc_hd__inv_2
XFILLER_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3500_ _3500_/A VGND VGND VPWR VPWR _3500_/Y sky130_fd_sc_hd__inv_2
X_4480_ _4480_/A _4480_/B VGND VGND VPWR VPWR _4481_/C sky130_fd_sc_hd__nand2_1
X_3431_ _3737_/A VGND VGND VPWR VPWR _3431_/X sky130_fd_sc_hd__clkbuf_2
X_3362_ _3370_/A VGND VGND VPWR VPWR _3737_/A sky130_fd_sc_hd__clkbuf_2
X_5101_ _3319_/X _5101_/D VGND VGND VPWR VPWR _5101_/Q sky130_fd_sc_hd__dfxtp_1
X_3293_ _3328_/A _3064_/X _3292_/Y VGND VGND VPWR VPWR _3294_/A sky130_fd_sc_hd__o21ai_1
X_5032_ _5047_/CLK _5032_/D VGND VGND VPWR VPWR _5032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4816_ _2444_/X _4816_/D VGND VGND VPWR VPWR _4816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4747_ _4634_/B _3041_/X _4715_/A _4745_/Y _4746_/X VGND VGND VPWR VPWR _4747_/X
+ sky130_fd_sc_hd__o221a_1
X_4678_ _4678_/A _4678_/B VGND VGND VPWR VPWR _4678_/X sky130_fd_sc_hd__or2_1
X_3629_ _4913_/Q VGND VGND VPWR VPWR _3630_/B sky130_fd_sc_hd__inv_2
Xoutput27 _4774_/Q VGND VGND VPWR VPWR DATA[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3980_ _3984_/A _3984_/B VGND VGND VPWR VPWR _3985_/B sky130_fd_sc_hd__or2_1
X_2931_ _5100_/Q _5137_/Q _2929_/Y _2930_/Y VGND VGND VPWR VPWR _3151_/A sky130_fd_sc_hd__o22a_1
X_2862_ _3488_/A _2861_/A _5062_/Q _2861_/Y VGND VGND VPWR VPWR _2922_/A sky130_fd_sc_hd__o22a_1
X_4601_ _4601_/A _4601_/B VGND VGND VPWR VPWR _4863_/D sky130_fd_sc_hd__nor2_1
X_2793_ _2703_/A _2774_/X _2775_/X VGND VGND VPWR VPWR _2795_/C sky130_fd_sc_hd__o21a_1
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A VGND VGND VPWR VPWR _4532_/Y sky130_fd_sc_hd__inv_2
X_4463_ _4611_/B _4856_/Q _4301_/Y _4610_/B _4857_/Q VGND VGND VPWR VPWR _4463_/X
+ sky130_fd_sc_hd__o32a_1
X_3414_ _3341_/A _3414_/A2 _3401_/X _3411_/Y VGND VGND VPWR VPWR _5083_/D sky130_fd_sc_hd__a211oi_1
X_4394_ _4793_/Q VGND VGND VPWR VPWR _4396_/A sky130_fd_sc_hd__inv_2
X_3345_ _3345_/A _3345_/B VGND VGND VPWR VPWR _3346_/B sky130_fd_sc_hd__or2_2
X_3276_ _3276_/A _3276_/B VGND VGND VPWR VPWR _3276_/Y sky130_fd_sc_hd__nand2_1
X_5015_ _5018_/CLK _5015_/D VGND VGND VPWR VPWR _5015_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3130_ _2986_/Y _3020_/X _3250_/A _3129_/X VGND VGND VPWR VPWR _3212_/A sky130_fd_sc_hd__o22a_2
XFILLER_67_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3061_ _3061_/A VGND VGND VPWR VPWR _3103_/A sky130_fd_sc_hd__inv_2
X_3963_ _3967_/A _3963_/B VGND VGND VPWR VPWR _3963_/X sky130_fd_sc_hd__or2_1
XFILLER_50_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3894_ _3985_/A _3894_/B _3894_/C VGND VGND VPWR VPWR _4969_/D sky130_fd_sc_hd__and3_1
X_2914_ _2914_/A _2914_/B _2914_/C VGND VGND VPWR VPWR _2914_/X sky130_fd_sc_hd__or3_1
X_2845_ _3523_/A _2845_/B VGND VGND VPWR VPWR _2846_/B sky130_fd_sc_hd__or2_1
X_2776_ _2691_/A _2774_/X _2775_/X VGND VGND VPWR VPWR _2780_/C sky130_fd_sc_hd__o21a_1
X_4515_ _4515_/A VGND VGND VPWR VPWR _4515_/Y sky130_fd_sc_hd__inv_2
X_4446_ _4446_/A _4446_/B VGND VGND VPWR VPWR _4450_/A sky130_fd_sc_hd__or2_1
X_4377_ _4569_/A _4564_/A VGND VGND VPWR VPWR _4387_/A sky130_fd_sc_hd__or2_1
X_3328_ _3328_/A _3328_/B VGND VGND VPWR VPWR _3329_/B sky130_fd_sc_hd__or2_1
X_3259_ _3259_/A _3259_/B VGND VGND VPWR VPWR _3259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2630_ _4939_/Q _2630_/B VGND VGND VPWR VPWR _2630_/Y sky130_fd_sc_hd__nor2_1
X_2561_ _4735_/A _3096_/B _4735_/C VGND VGND VPWR VPWR _2561_/X sky130_fd_sc_hd__o21a_1
X_4300_ _4857_/Q VGND VGND VPWR VPWR _4301_/B sky130_fd_sc_hd__inv_2
X_2492_ _4750_/X _4754_/Y VGND VGND VPWR VPWR _2492_/X sky130_fd_sc_hd__or2_1
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4231_ _4226_/A _4226_/B _4220_/X _4226_/Y VGND VGND VPWR VPWR _4914_/D sky130_fd_sc_hd__o211a_1
X_4162_ _4162_/A VGND VGND VPWR VPWR _4166_/A sky130_fd_sc_hd__inv_2
X_3113_ _3336_/A _3025_/X _3021_/Y _3337_/A _3112_/Y VGND VGND VPWR VPWR _3113_/X
+ sky130_fd_sc_hd__o32a_1
X_4093_ _4093_/A VGND VGND VPWR VPWR _4093_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3044_ _5111_/Q VGND VGND VPWR VPWR _3045_/A sky130_fd_sc_hd__inv_2
XFILLER_63_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4995_ _5028_/CLK _4995_/D VGND VGND VPWR VPWR _4995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3946_ _3786_/A _3945_/Y _3784_/A _3945_/A _3936_/X VGND VGND VPWR VPWR _4956_/D
+ sky130_fd_sc_hd__o221a_1
X_3877_ _3753_/Y _3893_/B _3893_/A _3876_/X VGND VGND VPWR VPWR _3887_/A sky130_fd_sc_hd__o31a_1
X_2828_ _4971_/Q _2781_/X _2796_/X VGND VGND VPWR VPWR _2830_/C sky130_fd_sc_hd__o21a_1
X_2759_ _2721_/A _2705_/X _2758_/X VGND VGND VPWR VPWR _2763_/A sky130_fd_sc_hd__o21a_1
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4429_ _4636_/B _4835_/Q _4637_/B _4834_/Q VGND VGND VPWR VPWR _4429_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_48_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4780_ _5139_/Q _4780_/D VGND VGND VPWR VPWR _4780_/Q sky130_fd_sc_hd__dfxtp_1
X_3800_ _4915_/Q _3799_/B _3799_/Y VGND VGND VPWR VPWR _3801_/A sky130_fd_sc_hd__a21oi_2
X_3731_ _4867_/Q VGND VGND VPWR VPWR _4091_/A sky130_fd_sc_hd__inv_2
X_3662_ _3668_/A _3662_/B VGND VGND VPWR VPWR _5009_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3593_ _3599_/A _3593_/B VGND VGND VPWR VPWR _5040_/D sky130_fd_sc_hd__nor2_1
X_2613_ _2756_/A _2613_/B VGND VGND VPWR VPWR _2613_/Y sky130_fd_sc_hd__nor2_1
X_2544_ _4720_/A _2539_/B _2517_/X _2539_/Y VGND VGND VPWR VPWR _4794_/D sky130_fd_sc_hd__o211a_1
X_2475_ _4684_/B _2475_/B VGND VGND VPWR VPWR _2475_/X sky130_fd_sc_hd__or2_1
X_4214_ _4210_/A _4210_/B _4177_/X _4210_/Y VGND VGND VPWR VPWR _4918_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4145_ _4014_/Y _4154_/B _4154_/A _4144_/X VGND VGND VPWR VPWR _4146_/A sky130_fd_sc_hd__o31a_1
XFILLER_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4076_ _3717_/B _4985_/Q _3717_/B _4985_/Q VGND VGND VPWR VPWR _4243_/A sky130_fd_sc_hd__a2bb2o_1
X_3027_ _3259_/A _3256_/A VGND VGND VPWR VPWR _3038_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4978_ _5018_/CLK _4978_/D VGND VGND VPWR VPWR _4978_/Q sky130_fd_sc_hd__dfxtp_2
X_3929_ _3609_/B _5033_/Q _3928_/Y VGND VGND VPWR VPWR _3930_/A sky130_fd_sc_hd__o21ai_1
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4901_ _5018_/CLK _4901_/D VGND VGND VPWR VPWR _4901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4832_ _5139_/Q _4832_/D VGND VGND VPWR VPWR _4832_/Q sky130_fd_sc_hd__dfxtp_1
X_4763_ _2755_/X _2746_/X _4770_/S VGND VGND VPWR VPWR _4780_/D sky130_fd_sc_hd__mux2_2
X_4694_ _4327_/X _2992_/X _4693_/X VGND VGND VPWR VPWR _4694_/Y sky130_fd_sc_hd__o21ai_1
X_3714_ _3714_/A _3714_/B VGND VGND VPWR VPWR _4986_/D sky130_fd_sc_hd__nor2_1
X_3645_ _3645_/A _3645_/B VGND VGND VPWR VPWR _5017_/D sky130_fd_sc_hd__nor2_1
X_3576_ _5048_/Q _3576_/B VGND VGND VPWR VPWR _5048_/D sky130_fd_sc_hd__nor2_1
X_2527_ _4709_/B _2521_/B _2517_/X _2521_/Y VGND VGND VPWR VPWR _4798_/D sky130_fd_sc_hd__o211a_1
X_2458_ _4618_/B _2981_/Y _2457_/X VGND VGND VPWR VPWR _2459_/A sky130_fd_sc_hd__o21ai_1
XFILLER_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2389_ _2389_/A VGND VGND VPWR VPWR _2391_/B sky130_fd_sc_hd__inv_2
X_4128_ _4886_/Q _4043_/B _4043_/Y VGND VGND VPWR VPWR _4129_/A sky130_fd_sc_hd__a21oi_2
X_4059_ _4131_/C _4059_/B VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__or2_1
XFILLER_56_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3430_ _3442_/A VGND VGND VPWR VPWR _3430_/X sky130_fd_sc_hd__buf_1
X_3361_ _3365_/A VGND VGND VPWR VPWR _3361_/X sky130_fd_sc_hd__buf_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5100_ _3322_/X _5100_/D VGND VGND VPWR VPWR _5100_/Q sky130_fd_sc_hd__dfxtp_1
X_3292_ _3292_/A _3292_/B VGND VGND VPWR VPWR _3292_/Y sky130_fd_sc_hd__nand2_1
X_5031_ _5047_/CLK _5031_/D VGND VGND VPWR VPWR _5031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4815_ _2446_/X _4815_/D VGND VGND VPWR VPWR _4815_/Q sky130_fd_sc_hd__dfxtp_1
X_4746_ _4634_/B _3041_/X _4635_/B _3045_/X VGND VGND VPWR VPWR _4746_/X sky130_fd_sc_hd__a211o_1
X_4677_ _4677_/A _4677_/B VGND VGND VPWR VPWR _4678_/B sky130_fd_sc_hd__or2_1
X_3628_ _3634_/A _3628_/B VGND VGND VPWR VPWR _5025_/D sky130_fd_sc_hd__nor2_1
Xoutput28 _4775_/Q VGND VGND VPWR VPWR DATA[3] sky130_fd_sc_hd__clkbuf_2
X_3559_ _3559_/A VGND VGND VPWR VPWR _3559_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2930_ _5137_/Q VGND VGND VPWR VPWR _2930_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2861_ _2861_/A VGND VGND VPWR VPWR _2861_/Y sky130_fd_sc_hd__inv_2
X_4600_ _4788_/Q _4414_/Y _4735_/A _4826_/Q VGND VGND VPWR VPWR _4601_/B sky130_fd_sc_hd__o22a_1
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2792_ _2666_/A _2791_/X _2772_/X VGND VGND VPWR VPWR _2795_/B sky130_fd_sc_hd__o21a_1
X_4531_ _4335_/A _4530_/Y _4331_/A _4530_/A _4501_/X VGND VGND VPWR VPWR _4884_/D
+ sky130_fd_sc_hd__o221a_1
X_4462_ _4819_/Q VGND VGND VPWR VPWR _4610_/B sky130_fd_sc_hd__inv_2
X_3413_ _3413_/A VGND VGND VPWR VPWR _3413_/X sky130_fd_sc_hd__buf_1
X_4393_ _4401_/A _4832_/Q _4401_/A _4832_/Q VGND VGND VPWR VPWR _4579_/A sky130_fd_sc_hd__a2bb2o_1
X_3344_ _3344_/A _3344_/B VGND VGND VPWR VPWR _3345_/B sky130_fd_sc_hd__or2_2
X_3275_ _3332_/A _3045_/X _3274_/Y VGND VGND VPWR VPWR _3276_/B sky130_fd_sc_hd__o21ai_1
X_5014_ _5018_/CLK _5014_/D VGND VGND VPWR VPWR _5014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4729_ _4791_/Q _5104_/Q VGND VGND VPWR VPWR _4729_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater36 _5028_/CLK VGND VGND VPWR VPWR _5047_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3060_ _5071_/Q _5108_/Q _3059_/Y VGND VGND VPWR VPWR _3061_/A sky130_fd_sc_hd__a21oi_2
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3962_ _3958_/A _3958_/B _3939_/X _3958_/Y VGND VGND VPWR VPWR _4951_/D sky130_fd_sc_hd__o211a_1
X_3893_ _3893_/A _3893_/B VGND VGND VPWR VPWR _3894_/C sky130_fd_sc_hd__nand2_1
X_2913_ _2910_/X _2912_/Y _2910_/X _2912_/Y VGND VGND VPWR VPWR _2914_/C sky130_fd_sc_hd__o2bb2a_1
X_2844_ input8/X input9/X VGND VGND VPWR VPWR _2845_/B sky130_fd_sc_hd__or2_1
X_4514_ _4618_/B _4850_/Q _4518_/B VGND VGND VPWR VPWR _4515_/A sky130_fd_sc_hd__o21ai_1
X_2775_ _2775_/A VGND VGND VPWR VPWR _2775_/X sky130_fd_sc_hd__clkbuf_2
X_4445_ _4445_/A _4542_/B VGND VGND VPWR VPWR _4446_/B sky130_fd_sc_hd__or2_1
X_4376_ _4431_/A _4836_/Q _4431_/A _4836_/Q VGND VGND VPWR VPWR _4564_/A sky130_fd_sc_hd__a2bb2o_1
X_3327_ _3327_/A _3327_/B VGND VGND VPWR VPWR _3328_/B sky130_fd_sc_hd__or2_1
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3258_ _3375_/A VGND VGND VPWR VPWR _3258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3189_ _3189_/A _3189_/B VGND VGND VPWR VPWR _3189_/X sky130_fd_sc_hd__or2_1
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2560_ _2560_/A VGND VGND VPWR VPWR _2560_/X sky130_fd_sc_hd__buf_1
X_2491_ _2497_/A VGND VGND VPWR VPWR _2491_/X sky130_fd_sc_hd__buf_1
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4230_ _4069_/A _4228_/Y _4067_/A _4228_/A _4229_/X VGND VGND VPWR VPWR _4915_/D
+ sky130_fd_sc_hd__o221a_1
X_4161_ _4481_/A _4161_/B _4161_/C VGND VGND VPWR VPWR _4932_/D sky130_fd_sc_hd__and3_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3112_ _5116_/Q VGND VGND VPWR VPWR _3112_/Y sky130_fd_sc_hd__inv_2
X_4092_ _4090_/A _4979_/Q _4090_/Y _4091_/Y VGND VGND VPWR VPWR _4093_/A sky130_fd_sc_hd__o2bb2a_1
X_3043_ _5074_/Q VGND VGND VPWR VPWR _3332_/A sky130_fd_sc_hd__clkinvlp_4
X_4994_ _5028_/CLK _4994_/D VGND VGND VPWR VPWR _4994_/Q sky130_fd_sc_hd__dfxtp_1
X_3945_ _3945_/A VGND VGND VPWR VPWR _3945_/Y sky130_fd_sc_hd__inv_2
X_3876_ _3586_/B _5043_/Q _3751_/Y _3584_/B _5044_/Q VGND VGND VPWR VPWR _3876_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2827_ _2827_/A _2827_/B _2827_/C _2827_/D VGND VGND VPWR VPWR _2830_/B sky130_fd_sc_hd__or4_4
X_2758_ _2758_/A VGND VGND VPWR VPWR _2758_/X sky130_fd_sc_hd__buf_1
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2689_ _2801_/A _2613_/B _2663_/X VGND VGND VPWR VPWR _2690_/D sky130_fd_sc_hd__o21a_1
X_4428_ _4428_/A VGND VGND VPWR VPWR _4634_/B sky130_fd_sc_hd__clkbuf_2
X_4359_ _4359_/A VGND VGND VPWR VPWR _4362_/A sky130_fd_sc_hd__inv_2
XFILLER_73_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3730_ _3736_/A _4090_/A VGND VGND VPWR VPWR _4979_/D sky130_fd_sc_hd__nor2_1
X_3661_ _4898_/Q VGND VGND VPWR VPWR _3662_/B sky130_fd_sc_hd__inv_2
X_3592_ _4929_/Q VGND VGND VPWR VPWR _3593_/B sky130_fd_sc_hd__inv_2
X_2612_ _2783_/A VGND VGND VPWR VPWR _2613_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2543_ _2543_/A VGND VGND VPWR VPWR _2543_/X sky130_fd_sc_hd__buf_1
XFILLER_5_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2474_ _2474_/A VGND VGND VPWR VPWR _2474_/X sky130_fd_sc_hd__buf_1
X_4213_ _4052_/A _4212_/Y _4050_/A _4212_/A _4190_/X VGND VGND VPWR VPWR _4919_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4144_ _3664_/B _5008_/Q _4012_/Y _3662_/B _5009_/Q VGND VGND VPWR VPWR _4144_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4075_ _4075_/A _4075_/B VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__or2_1
X_3026_ _3336_/A _3025_/X _5078_/Q _5115_/Q VGND VGND VPWR VPWR _3256_/A sky130_fd_sc_hd__o22a_1
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4977_ _5018_/CLK _4977_/D VGND VGND VPWR VPWR _4977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3928_ _3928_/A _3928_/B VGND VGND VPWR VPWR _3928_/Y sky130_fd_sc_hd__nand2_1
X_3859_ _3859_/A VGND VGND VPWR VPWR _3948_/B sky130_fd_sc_hd__inv_2
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4900_ _5018_/CLK _4900_/D VGND VGND VPWR VPWR _4900_/Q sky130_fd_sc_hd__dfxtp_1
X_4831_ _5139_/Q _4831_/D VGND VGND VPWR VPWR _4831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4762_ _2745_/X _2736_/X _4770_/S VGND VGND VPWR VPWR _4779_/D sky130_fd_sc_hd__mux2_2
XFILLER_33_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4693_ _4327_/X _2992_/X _4808_/Q _5121_/Q VGND VGND VPWR VPWR _4693_/X sky130_fd_sc_hd__a22o_1
X_3713_ _4875_/Q VGND VGND VPWR VPWR _3714_/B sky130_fd_sc_hd__inv_2
X_3644_ _4906_/Q VGND VGND VPWR VPWR _3645_/B sky130_fd_sc_hd__inv_2
X_3575_ _2899_/X _2900_/Y _5048_/Q _5049_/Q _3554_/X VGND VGND VPWR VPWR _5049_/D
+ sky130_fd_sc_hd__o221a_1
X_2526_ _2543_/A VGND VGND VPWR VPWR _2526_/X sky130_fd_sc_hd__buf_1
X_2457_ _2462_/A _4677_/B VGND VGND VPWR VPWR _2457_/X sky130_fd_sc_hd__or2_1
XFILLER_68_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2388_ _4811_/Q _5124_/Q _4679_/Y VGND VGND VPWR VPWR _2389_/A sky130_fd_sc_hd__a21oi_2
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4127_ _4127_/A _4127_/B VGND VGND VPWR VPWR _4131_/A sky130_fd_sc_hd__or2_1
XFILLER_56_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4058_ _3699_/B _4993_/Q _4127_/A _4056_/Y _4057_/X VGND VGND VPWR VPWR _4059_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3009_ _3340_/A _3008_/X _5082_/Q _5119_/Q VGND VGND VPWR VPWR _3235_/A sky130_fd_sc_hd__o22a_1
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3360_ _5100_/Q _3358_/Y _2929_/Y _3358_/A _3359_/X VGND VGND VPWR VPWR _5100_/D
+ sky130_fd_sc_hd__o221a_1
X_5030_ _5047_/CLK _5030_/D VGND VGND VPWR VPWR _5030_/Q sky130_fd_sc_hd__dfxtp_1
X_3291_ _3080_/A _3300_/B _3300_/A _3074_/A VGND VGND VPWR VPWR _3292_/B sky130_fd_sc_hd__a31o_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4814_ _2453_/X _4814_/D VGND VGND VPWR VPWR _4814_/Q sky130_fd_sc_hd__dfxtp_1
X_4745_ _4379_/X _3050_/X _4744_/X VGND VGND VPWR VPWR _4745_/Y sky130_fd_sc_hd__o21ai_1
X_4676_ _4676_/A VGND VGND VPWR VPWR _4677_/B sky130_fd_sc_hd__inv_2
X_3627_ _4914_/Q VGND VGND VPWR VPWR _3628_/B sky130_fd_sc_hd__inv_2
Xoutput29 _4776_/Q VGND VGND VPWR VPWR DATA[4] sky130_fd_sc_hd__clkbuf_2
X_3558_ _3558_/A VGND VGND VPWR VPWR _3558_/Y sky130_fd_sc_hd__inv_2
X_2509_ _2519_/A VGND VGND VPWR VPWR _2509_/X sky130_fd_sc_hd__buf_1
X_3489_ _3489_/A VGND VGND VPWR VPWR _3489_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2860_ input7/X _3494_/B _2922_/C VGND VGND VPWR VPWR _2861_/A sky130_fd_sc_hd__a21oi_2
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2791_ _2791_/A VGND VGND VPWR VPWR _2791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4530_ _4530_/A VGND VGND VPWR VPWR _4530_/Y sky130_fd_sc_hd__inv_2
X_4461_ _4461_/A VGND VGND VPWR VPWR _4611_/B sky130_fd_sc_hd__clkbuf_2
X_3412_ _5084_/Q _3411_/Y _3406_/X _3412_/C1 VGND VGND VPWR VPWR _5084_/D sky130_fd_sc_hd__o211a_1
X_4392_ _4794_/Q VGND VGND VPWR VPWR _4401_/A sky130_fd_sc_hd__inv_2
X_3343_ _3343_/A _3343_/B VGND VGND VPWR VPWR _3344_/B sky130_fd_sc_hd__or2_1
X_3274_ _3274_/A _3274_/B VGND VGND VPWR VPWR _3274_/Y sky130_fd_sc_hd__nand2_1
X_5013_ _5018_/CLK _5013_/D VGND VGND VPWR VPWR _5013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2989_ _5086_/Q VGND VGND VPWR VPWR _3344_/A sky130_fd_sc_hd__inv_1
X_4728_ _4728_/A _4728_/B VGND VGND VPWR VPWR _4740_/C sky130_fd_sc_hd__nand2_1
X_4659_ _4659_/A VGND VGND VPWR VPWR _4659_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater37 _5018_/CLK VGND VGND VPWR VPWR _5028_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3961_ _3803_/A _3960_/Y _3801_/A _3960_/A _3936_/X VGND VGND VPWR VPWR _4952_/D
+ sky130_fd_sc_hd__o221a_1
X_2912_ _2911_/Y _2907_/Y _2848_/B VGND VGND VPWR VPWR _2912_/Y sky130_fd_sc_hd__o21ai_1
X_3892_ _3753_/Y _3891_/Y _3753_/A _3891_/A _3359_/X VGND VGND VPWR VPWR _4970_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2843_ _5062_/Q VGND VGND VPWR VPWR _3488_/A sky130_fd_sc_hd__inv_2
X_2774_ _2774_/A VGND VGND VPWR VPWR _2774_/X sky130_fd_sc_hd__clkbuf_2
X_4513_ _4517_/A _4517_/B VGND VGND VPWR VPWR _4518_/B sky130_fd_sc_hd__or2_1
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4444_ _4444_/A VGND VGND VPWR VPWR _4542_/B sky130_fd_sc_hd__inv_2
X_4375_ _4798_/Q VGND VGND VPWR VPWR _4431_/A sky130_fd_sc_hd__inv_2
X_3326_ _3326_/A _3326_/B VGND VGND VPWR VPWR _3327_/B sky130_fd_sc_hd__or2_1
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3257_ _3336_/A _3025_/X _3256_/Y VGND VGND VPWR VPWR _3259_/B sky130_fd_sc_hd__o21ai_1
X_3188_ _3197_/A VGND VGND VPWR VPWR _3188_/X sky130_fd_sc_hd__buf_1
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2490_ _4687_/B _2484_/B _2486_/X _2484_/Y VGND VGND VPWR VPWR _4806_/D sky130_fd_sc_hd__o211a_1
X_4160_ _4160_/A _4160_/B VGND VGND VPWR VPWR _4161_/C sky130_fd_sc_hd__nand2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3111_ _5079_/Q VGND VGND VPWR VPWR _3337_/A sky130_fd_sc_hd__inv_2
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4091_ _4091_/A _4978_/Q VGND VGND VPWR VPWR _4091_/Y sky130_fd_sc_hd__nor2_4
X_3042_ _3333_/A _3041_/X _5075_/Q _5112_/Q VGND VGND VPWR VPWR _3276_/A sky130_fd_sc_hd__o22a_1
XFILLER_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4993_ _5028_/CLK _4993_/D VGND VGND VPWR VPWR _4993_/Q sky130_fd_sc_hd__dfxtp_1
X_3944_ _3618_/B _5029_/Q _3943_/Y VGND VGND VPWR VPWR _3945_/A sky130_fd_sc_hd__o21ai_1
X_3875_ _3766_/X _3775_/X _3923_/A _3874_/X VGND VGND VPWR VPWR _3893_/A sky130_fd_sc_hd__o31a_1
X_2826_ _4962_/Q _2777_/X _2778_/X VGND VGND VPWR VPWR _2827_/D sky130_fd_sc_hd__o21a_1
X_2757_ _2831_/A _2722_/X _2723_/X VGND VGND VPWR VPWR _2766_/A sky130_fd_sc_hd__o21a_1
X_2688_ _2831_/A _2606_/B _2659_/X VGND VGND VPWR VPWR _2690_/C sky130_fd_sc_hd__o21a_1
X_4427_ _4364_/X _4365_/Y _4426_/Y VGND VGND VPWR VPWR _4427_/Y sky130_fd_sc_hd__o21ai_1
X_4358_ _4803_/Q _4357_/B _4357_/Y VGND VGND VPWR VPWR _4359_/A sky130_fd_sc_hd__a21oi_2
XFILLER_48_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4289_ _4466_/A _4858_/Q _4466_/A _4858_/Q VGND VGND VPWR VPWR _4486_/B sky130_fd_sc_hd__a2bb2o_1
X_3309_ _3324_/D _3086_/X _3308_/X VGND VGND VPWR VPWR _3310_/A sky130_fd_sc_hd__o21ai_1
XFILLER_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3660_ _3660_/A _4899_/Q VGND VGND VPWR VPWR _5010_/D sky130_fd_sc_hd__and2_1
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3591_ _3599_/A _3591_/B VGND VGND VPWR VPWR _5041_/D sky130_fd_sc_hd__nor2_1
X_2611_ _2611_/A _2621_/B _2620_/D _2611_/D VGND VGND VPWR VPWR _2783_/A sky130_fd_sc_hd__nor4_2
X_2542_ _4740_/A _2541_/Y _4718_/A _2541_/A _2495_/X VGND VGND VPWR VPWR _4795_/D
+ sky130_fd_sc_hd__o221a_1
X_2473_ _2468_/A _2468_/B _2450_/X _2468_/Y VGND VGND VPWR VPWR _4810_/D sky130_fd_sc_hd__o211a_1
X_4212_ _4212_/A VGND VGND VPWR VPWR _4212_/Y sky130_fd_sc_hd__inv_2
X_4143_ _4019_/Y _4160_/B _4160_/A _4142_/X VGND VGND VPWR VPWR _4154_/A sky130_fd_sc_hd__o31a_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4074_ _4074_/A _4236_/A VGND VGND VPWR VPWR _4075_/B sky130_fd_sc_hd__or2_1
X_3025_ _3025_/A VGND VGND VPWR VPWR _3025_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4976_ _5018_/CLK _4976_/D VGND VGND VPWR VPWR _4976_/Q sky130_fd_sc_hd__dfxtp_1
X_3927_ _3865_/C _3933_/B _3795_/Y VGND VGND VPWR VPWR _3928_/B sky130_fd_sc_hd__o21ai_1
X_3858_ _3622_/B _5027_/Q _4916_/Q _3788_/Y VGND VGND VPWR VPWR _3859_/A sky130_fd_sc_hd__o22a_1
X_2809_ _4966_/Q _2783_/X _2798_/X VGND VGND VPWR VPWR _2810_/D sky130_fd_sc_hd__o21a_1
X_3789_ _4917_/Q _3787_/Y _4916_/Q _3788_/Y VGND VGND VPWR VPWR _3789_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4830_ _5139_/Q _4830_/D VGND VGND VPWR VPWR _4830_/Q sky130_fd_sc_hd__dfxtp_2
X_4761_ _2735_/X _2721_/X _4770_/S VGND VGND VPWR VPWR _4778_/D sky130_fd_sc_hd__mux2_2
XFILLER_60_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4692_ _4692_/A _4692_/B VGND VGND VPWR VPWR _4692_/X sky130_fd_sc_hd__or2_1
X_3712_ _3714_/A _3712_/B VGND VGND VPWR VPWR _4987_/D sky130_fd_sc_hd__nor2_1
X_3643_ _3645_/A _3643_/B VGND VGND VPWR VPWR _5018_/D sky130_fd_sc_hd__nor2_1
X_3574_ _3574_/A _3574_/B _3576_/B VGND VGND VPWR VPWR _5050_/D sky130_fd_sc_hd__nor3_1
X_2525_ _3384_/A VGND VGND VPWR VPWR _2543_/A sky130_fd_sc_hd__buf_1
X_2456_ _2474_/A VGND VGND VPWR VPWR _2456_/X sky130_fd_sc_hd__buf_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2387_ _4687_/Y _2387_/B VGND VGND VPWR VPWR _2391_/A sky130_fd_sc_hd__or2_1
X_4126_ _4126_/A _4215_/B VGND VGND VPWR VPWR _4127_/B sky130_fd_sc_hd__or2_1
XFILLER_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4057_ _3699_/B _4993_/Q _3701_/B _4992_/Q VGND VGND VPWR VPWR _4057_/X sky130_fd_sc_hd__a211o_1
X_3008_ _3008_/A VGND VGND VPWR VPWR _3008_/X sky130_fd_sc_hd__clkbuf_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4959_ _5018_/CLK _4959_/D VGND VGND VPWR VPWR _4959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3290_ _3290_/A VGND VGND VPWR VPWR _3300_/A sky130_fd_sc_hd__inv_2
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4813_ _2456_/X _4813_/D VGND VGND VPWR VPWR _4813_/Q sky130_fd_sc_hd__dfxtp_1
X_4744_ _4379_/X _3050_/X _4796_/Q _5109_/Q VGND VGND VPWR VPWR _4744_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4675_ _4317_/A _2981_/Y _4812_/Q _5125_/Q VGND VGND VPWR VPWR _4676_/A sky130_fd_sc_hd__o22a_1
X_3626_ _3634_/A _3626_/B VGND VGND VPWR VPWR _5026_/D sky130_fd_sc_hd__nor2_1
X_3557_ _3488_/A _3488_/B _3489_/Y _3576_/B VGND VGND VPWR VPWR _5062_/D sky130_fd_sc_hd__a211oi_1
Xoutput19 _4772_/Q VGND VGND VPWR VPWR DATA[0] sky130_fd_sc_hd__clkbuf_2
X_2508_ _4700_/A _2507_/B _2486_/X _2507_/Y VGND VGND VPWR VPWR _4803_/D sky130_fd_sc_hd__o211a_1
X_3488_ _3488_/A _3488_/B VGND VGND VPWR VPWR _3489_/A sky130_fd_sc_hd__or2_1
X_2439_ _2453_/A VGND VGND VPWR VPWR _2439_/X sky130_fd_sc_hd__buf_1
X_4109_ _3736_/B _4976_/Q _4099_/Y _3734_/B _4977_/Q VGND VGND VPWR VPWR _4109_/X
+ sky130_fd_sc_hd__o32a_1
X_5089_ _3394_/X _5089_/D VGND VGND VPWR VPWR _5089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2790_ _2746_/A _2770_/X _2758_/X VGND VGND VPWR VPWR _2795_/A sky130_fd_sc_hd__o21a_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4460_ _4614_/B _4853_/Q _4320_/A _4457_/Y _4459_/X VGND VGND VPWR VPWR _4460_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3411_ _3411_/A VGND VGND VPWR VPWR _3411_/Y sky130_fd_sc_hd__inv_2
X_4391_ _4391_/A VGND VGND VPWR VPWR _4424_/A sky130_fd_sc_hd__inv_2
X_3342_ _3342_/A _3342_/B VGND VGND VPWR VPWR _3343_/B sky130_fd_sc_hd__or2_1
X_3273_ _3286_/A _3058_/B _3108_/Y VGND VGND VPWR VPWR _3274_/B sky130_fd_sc_hd__o21ai_1
X_5012_ _5018_/CLK _5012_/D VGND VGND VPWR VPWR _5012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2988_ _5124_/Q VGND VGND VPWR VPWR _2988_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4727_ _4722_/A _4722_/B _4722_/Y VGND VGND VPWR VPWR _4728_/B sky130_fd_sc_hd__a21oi_4
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4658_ _4466_/A _2945_/A _4820_/Q _5133_/Q VGND VGND VPWR VPWR _4659_/A sky130_fd_sc_hd__o22a_1
X_3609_ _3611_/A _3609_/B VGND VGND VPWR VPWR _5033_/D sky130_fd_sc_hd__nor2_1
X_4589_ _4398_/Y _4588_/Y _4406_/A VGND VGND VPWR VPWR _4589_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater38 _5139_/Q VGND VGND VPWR VPWR _5018_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3960_ _3960_/A VGND VGND VPWR VPWR _3960_/Y sky130_fd_sc_hd__inv_2
X_2911_ _3516_/A VGND VGND VPWR VPWR _2911_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3891_ _3891_/A VGND VGND VPWR VPWR _3891_/Y sky130_fd_sc_hd__inv_2
X_2842_ _4771_/X VGND VGND VPWR VPWR _2842_/Y sky130_fd_sc_hd__inv_2
X_2773_ _2643_/A _2726_/X _2772_/X VGND VGND VPWR VPWR _2780_/B sky130_fd_sc_hd__o21a_1
X_4512_ _4507_/A _4507_/B _4264_/X _4507_/Y VGND VGND VPWR VPWR _4889_/D sky130_fd_sc_hd__o211a_1
X_4443_ _4628_/B _4842_/Q _4804_/Q _4345_/Y VGND VGND VPWR VPWR _4444_/A sky130_fd_sc_hd__o22a_1
X_4374_ _4428_/A _4837_/Q _4428_/A _4837_/Q VGND VGND VPWR VPWR _4569_/A sky130_fd_sc_hd__a2bb2o_1
X_3325_ _3325_/A _3461_/A VGND VGND VPWR VPWR _3326_/B sky130_fd_sc_hd__or2_2
X_3256_ _3256_/A _3256_/B VGND VGND VPWR VPWR _3256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3187_ _3180_/A _3180_/B _3186_/X _3180_/Y VGND VGND VPWR VPWR _5131_/D sky130_fd_sc_hd__o211a_1
XFILLER_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3110_ _3333_/A _3041_/X _3058_/A _3108_/Y _3109_/X VGND VGND VPWR VPWR _3110_/X
+ sky130_fd_sc_hd__o221a_1
X_4090_ _4090_/A _4979_/Q VGND VGND VPWR VPWR _4090_/Y sky130_fd_sc_hd__nor2_1
X_3041_ _3041_/A VGND VGND VPWR VPWR _3041_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4992_ _5028_/CLK _4992_/D VGND VGND VPWR VPWR _4992_/Q sky130_fd_sc_hd__dfxtp_1
X_3943_ _3943_/A _3943_/B VGND VGND VPWR VPWR _3943_/Y sky130_fd_sc_hd__nand2_1
X_3874_ _3766_/B _3868_/Y _3766_/X _3872_/X _3873_/X VGND VGND VPWR VPWR _3874_/X
+ sky130_fd_sc_hd__o221a_1
X_2825_ _2746_/A _2774_/X _2775_/X VGND VGND VPWR VPWR _2827_/C sky130_fd_sc_hd__o21a_1
XFILLER_31_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2756_ _2756_/A _2756_/B VGND VGND VPWR VPWR _2756_/X sky130_fd_sc_hd__or2_1
X_2687_ _4960_/Q VGND VGND VPWR VPWR _2831_/A sky130_fd_sc_hd__clkbuf_2
X_4426_ _4631_/B _4839_/Q _4632_/B _4838_/Q VGND VGND VPWR VPWR _4426_/Y sky130_fd_sc_hd__o22ai_1
X_4357_ _4803_/Q _4357_/B VGND VGND VPWR VPWR _4357_/Y sky130_fd_sc_hd__nor2_1
X_3308_ _3308_/A _3308_/B VGND VGND VPWR VPWR _3308_/X sky130_fd_sc_hd__or2_1
X_4288_ _4820_/Q VGND VGND VPWR VPWR _4466_/A sky130_fd_sc_hd__inv_2
X_3239_ _3241_/A VGND VGND VPWR VPWR _3239_/X sky130_fd_sc_hd__buf_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3590_ _4930_/Q VGND VGND VPWR VPWR _3591_/B sky130_fd_sc_hd__inv_2
X_2610_ _2610_/A _4968_/Q _2621_/C _4970_/Q VGND VGND VPWR VPWR _2611_/D sky130_fd_sc_hd__or4b_4
X_2541_ _2541_/A VGND VGND VPWR VPWR _2541_/Y sky130_fd_sc_hd__inv_2
X_2472_ _2474_/A VGND VGND VPWR VPWR _2472_/X sky130_fd_sc_hd__buf_1
XFILLER_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4211_ _3701_/B _4992_/Q _4210_/Y VGND VGND VPWR VPWR _4212_/A sky130_fd_sc_hd__o21ai_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4142_ _3668_/B _5006_/Q _4017_/Y _3666_/B _5007_/Q VGND VGND VPWR VPWR _4142_/X
+ sky130_fd_sc_hd__o32a_1
X_4073_ _3714_/B _4986_/Q _3714_/B _4986_/Q VGND VGND VPWR VPWR _4236_/A sky130_fd_sc_hd__a2bb2o_1
X_3024_ _5115_/Q VGND VGND VPWR VPWR _3025_/A sky130_fd_sc_hd__inv_2
XFILLER_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4975_ _5018_/CLK _4975_/D VGND VGND VPWR VPWR _4975_/Q sky130_fd_sc_hd__dfxtp_1
X_3926_ _3926_/A VGND VGND VPWR VPWR _3933_/B sky130_fd_sc_hd__inv_2
XFILLER_50_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3857_ _3857_/A VGND VGND VPWR VPWR _3860_/A sky130_fd_sc_hd__inv_2
X_2808_ _4969_/Q _2781_/X _2796_/X VGND VGND VPWR VPWR _2810_/C sky130_fd_sc_hd__o21a_1
X_3788_ _5027_/Q VGND VGND VPWR VPWR _3788_/Y sky130_fd_sc_hd__inv_2
X_2739_ _4943_/Q _2726_/X _2707_/X VGND VGND VPWR VPWR _2742_/B sky130_fd_sc_hd__o21a_1
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4409_ _4791_/Q _4408_/B _4408_/Y VGND VGND VPWR VPWR _4410_/A sky130_fd_sc_hd__a21oi_2
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4760_ _2720_/X _2703_/X _4770_/S VGND VGND VPWR VPWR _4777_/D sky130_fd_sc_hd__mux2_2
X_4691_ _4624_/B _3004_/X _4687_/Y _4689_/Y _4690_/X VGND VGND VPWR VPWR _4692_/B
+ sky130_fd_sc_hd__o221a_1
X_3711_ _4876_/Q VGND VGND VPWR VPWR _3712_/B sky130_fd_sc_hd__inv_2
X_3642_ _4907_/Q VGND VGND VPWR VPWR _3643_/B sky130_fd_sc_hd__inv_2
X_3573_ _2899_/X _2900_/Y _2895_/Y VGND VGND VPWR VPWR _3574_/B sky130_fd_sc_hd__o21a_1
X_2524_ _4709_/A _2523_/B _2517_/X _2523_/Y VGND VGND VPWR VPWR _4799_/D sky130_fd_sc_hd__o211a_1
X_2455_ _3459_/A VGND VGND VPWR VPWR _2474_/A sky130_fd_sc_hd__buf_1
X_2386_ _4752_/Y _4754_/Y VGND VGND VPWR VPWR _2387_/B sky130_fd_sc_hd__or2_1
X_4125_ _4125_/A VGND VGND VPWR VPWR _4215_/B sky130_fd_sc_hd__inv_2
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4056_ _4880_/Q _4053_/Y _4055_/X VGND VGND VPWR VPWR _4056_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3007_ _5119_/Q VGND VGND VPWR VPWR _3008_/A sky130_fd_sc_hd__inv_2
XFILLER_36_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4958_ _5018_/CLK _4958_/D VGND VGND VPWR VPWR _4958_/Q sky130_fd_sc_hd__dfxtp_1
X_3909_ _3909_/A VGND VGND VPWR VPWR _3909_/Y sky130_fd_sc_hd__inv_2
X_4889_ _5047_/CLK _4889_/D VGND VGND VPWR VPWR _4889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4812_ _2461_/X _4812_/D VGND VGND VPWR VPWR _4812_/Q sky130_fd_sc_hd__dfxtp_1
X_4743_ _4364_/X _3030_/X _4742_/X VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__o21ai_1
X_4674_ _4674_/A VGND VGND VPWR VPWR _4677_/A sky130_fd_sc_hd__inv_2
X_3625_ _4915_/Q VGND VGND VPWR VPWR _3626_/B sky130_fd_sc_hd__inv_2
X_3556_ _3556_/A VGND VGND VPWR VPWR _3576_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2507_ _4700_/A _2507_/B VGND VGND VPWR VPWR _2507_/Y sky130_fd_sc_hd__nand2_1
X_3487_ _3487_/A _3558_/A VGND VGND VPWR VPWR _3488_/B sky130_fd_sc_hd__or2_1
X_2438_ _4668_/A _2432_/B _2417_/X _2432_/Y VGND VGND VPWR VPWR _4818_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5088_ _3396_/X _5088_/D VGND VGND VPWR VPWR _5088_/Q sky130_fd_sc_hd__dfxtp_1
X_4108_ _4108_/A VGND VGND VPWR VPWR _4266_/A sky130_fd_sc_hd__inv_2
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4039_ _3687_/B _4998_/Q _3687_/B _4998_/Q VGND VGND VPWR VPWR _4192_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3410_ _3413_/A VGND VGND VPWR VPWR _3410_/X sky130_fd_sc_hd__buf_1
X_4390_ _4795_/Q _4389_/B _4389_/Y VGND VGND VPWR VPWR _4391_/A sky130_fd_sc_hd__a21oi_2
X_3341_ _3341_/A _3341_/B VGND VGND VPWR VPWR _3342_/B sky130_fd_sc_hd__or2_1
X_3272_ _3289_/A VGND VGND VPWR VPWR _3272_/X sky130_fd_sc_hd__buf_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5011_ _5018_/CLK _5011_/D VGND VGND VPWR VPWR _5011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2987_ _5087_/Q VGND VGND VPWR VPWR _3345_/A sky130_fd_sc_hd__clkinv_1
X_4726_ _4721_/A _4721_/B _4721_/Y VGND VGND VPWR VPWR _4728_/A sky130_fd_sc_hd__a21oi_4
X_4657_ _4657_/A VGND VGND VPWR VPWR _4657_/Y sky130_fd_sc_hd__inv_2
X_3608_ _3608_/A VGND VGND VPWR VPWR _3609_/B sky130_fd_sc_hd__buf_1
X_4588_ _4588_/A VGND VGND VPWR VPWR _4588_/Y sky130_fd_sc_hd__inv_2
X_3539_ _3479_/A _3538_/X _3479_/A _3538_/X VGND VGND VPWR VPWR _3542_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2910_ _5052_/Q VGND VGND VPWR VPWR _2910_/X sky130_fd_sc_hd__buf_1
XFILLER_16_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3890_ _3586_/B _5043_/Q _3894_/B VGND VGND VPWR VPWR _3891_/A sky130_fd_sc_hd__o21ai_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2841_ _5139_/Q _3318_/C _3554_/X _2923_/B VGND VGND VPWR VPWR _5139_/D sky130_fd_sc_hd__a31o_1
XFILLER_31_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2772_ _2772_/A VGND VGND VPWR VPWR _2772_/X sky130_fd_sc_hd__buf_1
X_4511_ _4510_/A _4509_/Y _4510_/Y _4509_/A _4501_/X VGND VGND VPWR VPWR _4890_/D
+ sky130_fd_sc_hd__o221a_1
X_4442_ _4804_/Q VGND VGND VPWR VPWR _4628_/B sky130_fd_sc_hd__inv_2
X_4373_ _4799_/Q VGND VGND VPWR VPWR _4428_/A sky130_fd_sc_hd__inv_2
X_3324_ _3324_/A _3324_/B _3324_/C _3324_/D VGND VGND VPWR VPWR _3461_/A sky130_fd_sc_hd__or4_4
X_3255_ _3038_/B _3264_/B _3106_/Y VGND VGND VPWR VPWR _3256_/B sky130_fd_sc_hd__o21ai_1
X_3186_ _3375_/A VGND VGND VPWR VPWR _3186_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4709_ _4709_/A _4709_/B VGND VGND VPWR VPWR _4715_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3040_ _5112_/Q VGND VGND VPWR VPWR _3041_/A sky130_fd_sc_hd__inv_2
XFILLER_75_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4991_ _5028_/CLK _4991_/D VGND VGND VPWR VPWR _4991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3942_ _3952_/A _3861_/B _3790_/Y VGND VGND VPWR VPWR _3943_/B sky130_fd_sc_hd__o21ai_1
X_3873_ _3591_/B _5041_/Q _3762_/Y _3588_/B _5042_/Q VGND VGND VPWR VPWR _3873_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2824_ _2703_/A _2791_/X _2772_/X VGND VGND VPWR VPWR _2827_/B sky130_fd_sc_hd__o21a_1
X_2755_ _2755_/A _2755_/B _2755_/C _2755_/D VGND VGND VPWR VPWR _2755_/X sky130_fd_sc_hd__or4_4
XFILLER_8_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2686_ _2686_/A _2686_/B _2686_/C _2686_/D VGND VGND VPWR VPWR _2690_/B sky130_fd_sc_hd__or4_4
X_4425_ _4424_/A _4579_/A _4400_/Y _4403_/X _4424_/X VGND VGND VPWR VPWR _4577_/A
+ sky130_fd_sc_hd__o311a_2
X_4356_ _4841_/Q VGND VGND VPWR VPWR _4357_/B sky130_fd_sc_hd__inv_2
X_3307_ _3312_/A VGND VGND VPWR VPWR _3307_/X sky130_fd_sc_hd__buf_1
XFILLER_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4287_ _4287_/A VGND VGND VPWR VPWR _4287_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3238_ _3237_/A _3237_/B _3223_/X _3237_/Y VGND VGND VPWR VPWR _5120_/D sky130_fd_sc_hd__o211a_1
X_3169_ _3354_/A _2945_/X _3168_/X VGND VGND VPWR VPWR _3170_/A sky130_fd_sc_hd__o21ai_1
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2540_ _4640_/B _3064_/X _2539_/Y VGND VGND VPWR VPWR _2541_/A sky130_fd_sc_hd__o21ai_1
X_2471_ _2391_/B _2470_/Y _2389_/A _2470_/A _2423_/X VGND VGND VPWR VPWR _4811_/D
+ sky130_fd_sc_hd__o221a_1
X_4210_ _4210_/A _4210_/B VGND VGND VPWR VPWR _4210_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4141_ _4032_/X _4041_/X _4192_/A _4140_/X VGND VGND VPWR VPWR _4160_/A sky130_fd_sc_hd__o31a_1
XFILLER_68_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4072_ _4072_/A VGND VGND VPWR VPWR _4074_/A sky130_fd_sc_hd__inv_2
X_3023_ _5078_/Q VGND VGND VPWR VPWR _3336_/A sky130_fd_sc_hd__clkinvlp_4
XFILLER_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4974_ _5018_/CLK _4974_/D VGND VGND VPWR VPWR _4974_/Q sky130_fd_sc_hd__dfxtp_1
X_3925_ _3952_/A _3865_/A _3793_/B VGND VGND VPWR VPWR _3926_/A sky130_fd_sc_hd__o21ai_1
X_3856_ _4917_/Q _3787_/Y _3620_/B _5028_/Q VGND VGND VPWR VPWR _3857_/A sky130_fd_sc_hd__o22a_1
X_2807_ _2807_/A _2807_/B _2807_/C _2807_/D VGND VGND VPWR VPWR _2810_/B sky130_fd_sc_hd__or4_4
X_3787_ _5028_/Q VGND VGND VPWR VPWR _3787_/Y sky130_fd_sc_hd__inv_2
X_2738_ _2691_/A _2705_/X _2693_/X VGND VGND VPWR VPWR _2742_/A sky130_fd_sc_hd__o21a_1
X_4408_ _4791_/Q _4408_/B VGND VGND VPWR VPWR _4408_/Y sky130_fd_sc_hd__nor2_1
X_2669_ _4944_/Q _2638_/X _2590_/A VGND VGND VPWR VPWR _2674_/A sky130_fd_sc_hd__o21a_1
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4339_ _4339_/A VGND VGND VPWR VPWR _4342_/A sky130_fd_sc_hd__inv_2
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3710_ _3714_/A _3710_/B VGND VGND VPWR VPWR _4988_/D sky130_fd_sc_hd__nor2_1
X_4690_ _4624_/B _3004_/X _4625_/B _3008_/X VGND VGND VPWR VPWR _4690_/X sky130_fd_sc_hd__a211o_1
X_3641_ _3645_/A _3641_/B VGND VGND VPWR VPWR _5019_/D sky130_fd_sc_hd__nor2_1
X_3572_ _3525_/A _3574_/A _3476_/A _3554_/X VGND VGND VPWR VPWR _5051_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2523_ _4709_/A _2523_/B VGND VGND VPWR VPWR _2523_/Y sky130_fd_sc_hd__nand2_1
X_2454_ _4672_/B _2448_/B _2450_/X _2448_/Y VGND VGND VPWR VPWR _4814_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4124_ _3706_/B _4990_/Q _4879_/Q _4054_/Y VGND VGND VPWR VPWR _4125_/A sky130_fd_sc_hd__o22a_1
Xinput1 dec_rate[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4055_ _4880_/Q _4053_/Y _4879_/Q _4054_/Y VGND VGND VPWR VPWR _4055_/X sky130_fd_sc_hd__a22o_1
X_3006_ _5082_/Q VGND VGND VPWR VPWR _3340_/A sky130_fd_sc_hd__clkinvlp_4
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4957_ _5018_/CLK _4957_/D VGND VGND VPWR VPWR _4957_/Q sky130_fd_sc_hd__dfxtp_1
X_3908_ _3759_/B _3907_/Y _3758_/A _3907_/A _3902_/X VGND VGND VPWR VPWR _4966_/D
+ sky130_fd_sc_hd__o221a_1
X_4888_ _5047_/CLK _4888_/D VGND VGND VPWR VPWR _4888_/Q sky130_fd_sc_hd__dfxtp_1
X_3839_ _3656_/B _5012_/Q _4901_/Q _3838_/Y VGND VGND VPWR VPWR _3839_/X sky130_fd_sc_hd__o22a_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4811_ _2464_/X _4811_/D VGND VGND VPWR VPWR _4811_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4742_ _4364_/X _3030_/X _4800_/Q _5113_/Q VGND VGND VPWR VPWR _4742_/X sky130_fd_sc_hd__a22o_1
X_4673_ _4617_/B _2976_/Y _4312_/X _5126_/Q VGND VGND VPWR VPWR _4674_/A sky130_fd_sc_hd__o22a_1
X_3624_ _3669_/A VGND VGND VPWR VPWR _3634_/A sky130_fd_sc_hd__clkbuf_2
X_3555_ _5063_/Q _3489_/Y _2880_/Y _3489_/A _3554_/X VGND VGND VPWR VPWR _5063_/D
+ sky130_fd_sc_hd__o221a_1
X_3486_ _3486_/A _3486_/B VGND VGND VPWR VPWR _3558_/A sky130_fd_sc_hd__or2_1
X_2506_ _4630_/B _3025_/X _2505_/Y VGND VGND VPWR VPWR _2507_/B sky130_fd_sc_hd__o21ai_1
X_2437_ _2453_/A VGND VGND VPWR VPWR _2437_/X sky130_fd_sc_hd__buf_1
X_5087_ _3400_/X _5087_/D VGND VGND VPWR VPWR _5087_/Q sky130_fd_sc_hd__dfxtp_1
X_4107_ _3740_/B _4975_/Q _4106_/Y VGND VGND VPWR VPWR _4108_/A sky130_fd_sc_hd__o21ai_2
X_4038_ _4038_/A VGND VGND VPWR VPWR _4040_/A sky130_fd_sc_hd__inv_2
XFILLER_52_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3340_ _3340_/A _3340_/B VGND VGND VPWR VPWR _3341_/B sky130_fd_sc_hd__or2_1
X_5010_ _5047_/CLK _5010_/D VGND VGND VPWR VPWR _5010_/Q sky130_fd_sc_hd__dfxtp_1
X_3271_ _3368_/A VGND VGND VPWR VPWR _3289_/A sky130_fd_sc_hd__buf_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2986_ _5087_/Q _5124_/Q VGND VGND VPWR VPWR _2986_/Y sky130_fd_sc_hd__nor2_2
X_4725_ _4640_/B _3064_/X _4716_/Y _4638_/B _3076_/Y VGND VGND VPWR VPWR _4725_/X
+ sky130_fd_sc_hd__o32a_1
X_4656_ _4821_/Q _5134_/Q _4655_/Y VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__a21oi_2
X_4587_ _4587_/A _4587_/B VGND VGND VPWR VPWR _4588_/A sky130_fd_sc_hd__nand2_1
X_3607_ _4922_/Q VGND VGND VPWR VPWR _3608_/A sky130_fd_sc_hd__inv_2
X_3538_ _3517_/A _3517_/B _3517_/X VGND VGND VPWR VPWR _3538_/X sky130_fd_sc_hd__a21bo_1
X_3469_ _3320_/X _3469_/A2 _3090_/X _4578_/A _3468_/Y VGND VGND VPWR VPWR _5065_/D
+ sky130_fd_sc_hd__o311a_1
X_5139_ _5139_/CLK _5139_/D VGND VGND VPWR VPWR _5139_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2840_ _2840_/A _2840_/B _2840_/C _2840_/D VGND VGND VPWR VPWR _2840_/X sky130_fd_sc_hd__or4_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _2736_/A _2770_/X _2758_/X VGND VGND VPWR VPWR _2780_/A sky130_fd_sc_hd__o21a_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4510_ _4510_/A VGND VGND VPWR VPWR _4510_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4441_ _4441_/A VGND VGND VPWR VPWR _4445_/A sky130_fd_sc_hd__inv_2
X_4372_ _4372_/A _4372_/B VGND VGND VPWR VPWR _4372_/X sky130_fd_sc_hd__or2_1
X_3323_ _3323_/A VGND VGND VPWR VPWR _3324_/B sky130_fd_sc_hd__inv_1
X_3254_ _3254_/A VGND VGND VPWR VPWR _3264_/B sky130_fd_sc_hd__inv_2
X_3185_ _4176_/A VGND VGND VPWR VPWR _3375_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2969_ _3349_/A _2968_/X _5091_/Q _5128_/Q VGND VGND VPWR VPWR _3201_/A sky130_fd_sc_hd__o22a_1
X_4708_ _4431_/A _3045_/A _4798_/Q _5111_/Q VGND VGND VPWR VPWR _4709_/B sky130_fd_sc_hd__o22a_1
X_4639_ _4639_/A VGND VGND VPWR VPWR _4644_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4990_ _5028_/CLK _4990_/D VGND VGND VPWR VPWR _4990_/Q sky130_fd_sc_hd__dfxtp_1
X_3941_ _3941_/A VGND VGND VPWR VPWR _3943_/A sky130_fd_sc_hd__inv_2
X_3872_ _3597_/B _5038_/Q _3775_/A _3870_/Y _3871_/X VGND VGND VPWR VPWR _3872_/X
+ sky130_fd_sc_hd__o221a_1
X_2823_ _2786_/A _2770_/X _2758_/A VGND VGND VPWR VPWR _2827_/A sky130_fd_sc_hd__o21a_1
X_2754_ _4962_/Q _2718_/X _2733_/X VGND VGND VPWR VPWR _2755_/D sky130_fd_sc_hd__o21a_1
X_2685_ _2721_/A _2624_/B _2590_/D VGND VGND VPWR VPWR _2686_/D sky130_fd_sc_hd__o21a_1
X_4424_ _4424_/A _4579_/A _4424_/C _4580_/A VGND VGND VPWR VPWR _4424_/X sky130_fd_sc_hd__or4_4
X_4355_ _4619_/B _4849_/Q _4620_/B _4848_/Q _4354_/X VGND VGND VPWR VPWR _4355_/X
+ sky130_fd_sc_hd__o221a_1
X_3306_ _3300_/A _3300_/B _3287_/X _3301_/A VGND VGND VPWR VPWR _5105_/D sky130_fd_sc_hd__o211a_1
X_4286_ _4821_/Q _4285_/B _4285_/Y VGND VGND VPWR VPWR _4287_/A sky130_fd_sc_hd__a21oi_2
X_3237_ _3237_/A _3237_/B VGND VGND VPWR VPWR _3237_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3168_ _3173_/A _3168_/B VGND VGND VPWR VPWR _3168_/X sky130_fd_sc_hd__or2_1
X_3099_ _5067_/Q VGND VGND VPWR VPWR _3325_/A sky130_fd_sc_hd__clkinvlp_2
XFILLER_80_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2470_ _2470_/A VGND VGND VPWR VPWR _2470_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4140_ _4032_/B _4134_/Y _4032_/X _4138_/X _4139_/X VGND VGND VPWR VPWR _4140_/X
+ sky130_fd_sc_hd__o221a_1
X_4071_ _3712_/B _4987_/Q _4876_/Q _4070_/Y VGND VGND VPWR VPWR _4072_/A sky130_fd_sc_hd__o22a_1
X_3022_ _5079_/Q _5116_/Q _3021_/Y VGND VGND VPWR VPWR _3259_/A sky130_fd_sc_hd__a21oi_2
XFILLER_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4973_ _5018_/CLK _4973_/D VGND VGND VPWR VPWR _4973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3924_ _3985_/A _3924_/B _3924_/C VGND VGND VPWR VPWR _4961_/D sky130_fd_sc_hd__and3_1
XFILLER_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3855_ _3809_/X _3818_/X _3984_/A _3854_/X VGND VGND VPWR VPWR _3952_/A sky130_fd_sc_hd__o31a_2
X_2806_ _2831_/A _2777_/X _2778_/X VGND VGND VPWR VPWR _2807_/D sky130_fd_sc_hd__o21a_1
X_3786_ _3786_/A _3941_/A VGND VGND VPWR VPWR _3861_/A sky130_fd_sc_hd__or2_1
X_2737_ _2811_/A _2722_/X _2723_/X VGND VGND VPWR VPWR _2745_/A sky130_fd_sc_hd__o21a_1
X_2668_ _2746_/A _2645_/X _2647_/X VGND VGND VPWR VPWR _2679_/A sky130_fd_sc_hd__o21a_1
X_4407_ _4829_/Q VGND VGND VPWR VPWR _4408_/B sky130_fd_sc_hd__inv_2
X_2599_ _4972_/Q _4971_/Q _4973_/Q VGND VGND VPWR VPWR _2600_/C sky130_fd_sc_hd__or3b_2
X_4338_ _4337_/A _4845_/Q _4337_/A _4845_/Q VGND VGND VPWR VPWR _4339_/A sky130_fd_sc_hd__o2bb2a_1
X_4269_ _4269_/A VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3640_ _4908_/Q VGND VGND VPWR VPWR _3641_/B sky130_fd_sc_hd__inv_2
X_3571_ _2910_/X _3477_/B _3478_/B _3554_/X VGND VGND VPWR VPWR _5052_/D sky130_fd_sc_hd__o211a_1
X_2522_ _4635_/B _3045_/X _2521_/Y VGND VGND VPWR VPWR _2523_/B sky130_fd_sc_hd__o21ai_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2453_ _2453_/A VGND VGND VPWR VPWR _2453_/X sky130_fd_sc_hd__buf_1
X_4123_ _4123_/A VGND VGND VPWR VPWR _4126_/A sky130_fd_sc_hd__inv_2
Xinput2 dec_rate[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4054_ _4990_/Q VGND VGND VPWR VPWR _4054_/Y sky130_fd_sc_hd__inv_2
X_3005_ _5083_/Q _5120_/Q _3341_/A _3004_/X VGND VGND VPWR VPWR _3237_/A sky130_fd_sc_hd__o22a_1
XFILLER_64_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4956_ _5018_/CLK _4956_/D VGND VGND VPWR VPWR _4956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3907_ _3907_/A VGND VGND VPWR VPWR _3907_/Y sky130_fd_sc_hd__inv_2
X_4887_ _5047_/CLK _4887_/D VGND VGND VPWR VPWR _4887_/Q sky130_fd_sc_hd__dfxtp_1
X_3838_ _5012_/Q VGND VGND VPWR VPWR _3838_/Y sky130_fd_sc_hd__inv_2
X_3769_ _3916_/A _3911_/A VGND VGND VPWR VPWR _3775_/A sky130_fd_sc_hd__or2_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ _2472_/X _4810_/D VGND VGND VPWR VPWR _4810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4741_ _4740_/A _4740_/B _4724_/Y _4725_/X _4740_/X VGND VGND VPWR VPWR _4741_/X
+ sky130_fd_sc_hd__o311a_2
X_4672_ _4672_/A _4672_/B VGND VGND VPWR VPWR _4678_/A sky130_fd_sc_hd__nand2_1
X_3623_ _3737_/A VGND VGND VPWR VPWR _3669_/A sky130_fd_sc_hd__buf_2
X_3554_ _3559_/A VGND VGND VPWR VPWR _3554_/X sky130_fd_sc_hd__clkbuf_2
X_2505_ _4700_/B _2505_/B VGND VGND VPWR VPWR _2505_/Y sky130_fd_sc_hd__nand2_1
X_3485_ _3485_/A _3562_/A VGND VGND VPWR VPWR _3486_/B sky130_fd_sc_hd__or2_1
X_2436_ _3459_/A VGND VGND VPWR VPWR _2453_/A sky130_fd_sc_hd__buf_1
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5086_ _3403_/X _5086_/D VGND VGND VPWR VPWR _5086_/Q sky130_fd_sc_hd__dfxtp_1
X_4106_ _4863_/Q _4103_/Y _4105_/X VGND VGND VPWR VPWR _4106_/Y sky130_fd_sc_hd__o21ai_1
X_4037_ _3685_/B _4999_/Q _4888_/Q _4036_/Y VGND VGND VPWR VPWR _4038_/A sky130_fd_sc_hd__o22a_1
XFILLER_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4939_ _5018_/CLK _4939_/D VGND VGND VPWR VPWR _4939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3270_ _3036_/A _3254_/A _3258_/X _3264_/X VGND VGND VPWR VPWR _5113_/D sky130_fd_sc_hd__o211a_1
XFILLER_78_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4724_ _4724_/A VGND VGND VPWR VPWR _4724_/Y sky130_fd_sc_hd__inv_2
X_2985_ _2985_/A _2985_/B VGND VGND VPWR VPWR _2985_/X sky130_fd_sc_hd__or2_1
X_4655_ _4821_/Q _5134_/Q VGND VGND VPWR VPWR _4655_/Y sky130_fd_sc_hd__nor2_1
X_3606_ _3611_/A _3606_/B VGND VGND VPWR VPWR _5034_/D sky130_fd_sc_hd__nor2_1
X_4586_ _4582_/A _4582_/B _4562_/X _4582_/Y VGND VGND VPWR VPWR _4869_/D sky130_fd_sc_hd__o211a_1
X_3537_ _5053_/Q _3536_/Y _5053_/Q _3536_/Y VGND VGND VPWR VPWR _3542_/B sky130_fd_sc_hd__a2bb2o_1
X_3468_ _3320_/X _3468_/A2 _3090_/X VGND VGND VPWR VPWR _3468_/Y sky130_fd_sc_hd__o21ai_1
X_3399_ _3444_/A VGND VGND VPWR VPWR _3413_/A sky130_fd_sc_hd__buf_1
X_2419_ _2428_/A VGND VGND VPWR VPWR _2419_/X sky130_fd_sc_hd__buf_1
X_5138_ _5139_/CLK _5138_/D VGND VGND VPWR VPWR _5138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5069_ _3453_/X _5069_/D VGND VGND VPWR VPWR _5069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _2770_/A VGND VGND VPWR VPWR _2770_/X sky130_fd_sc_hd__clkbuf_2
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4440_ _4343_/X _4344_/Y _4626_/B _4843_/Q VGND VGND VPWR VPWR _4441_/A sky130_fd_sc_hd__o22a_1
X_4371_ _4371_/A _4561_/A VGND VGND VPWR VPWR _4372_/B sky130_fd_sc_hd__or2_1
X_3322_ _3365_/A VGND VGND VPWR VPWR _3322_/X sky130_fd_sc_hd__buf_1
X_3253_ _3286_/A _3058_/X _3110_/X VGND VGND VPWR VPWR _3254_/A sky130_fd_sc_hd__o21ai_1
X_3184_ _3197_/A VGND VGND VPWR VPWR _3184_/X sky130_fd_sc_hd__buf_1
XFILLER_66_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2968_ _2968_/A VGND VGND VPWR VPWR _2968_/X sky130_fd_sc_hd__clkbuf_2
X_4707_ _4428_/A _3041_/A _4799_/Q _5112_/Q VGND VGND VPWR VPWR _4709_/A sky130_fd_sc_hd__o22a_1
X_2899_ _2903_/A VGND VGND VPWR VPWR _2899_/X sky130_fd_sc_hd__buf_1
X_4638_ _4638_/A _4638_/B VGND VGND VPWR VPWR _4833_/D sky130_fd_sc_hd__nor2_1
X_4569_ _4569_/A VGND VGND VPWR VPWR _4569_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3940_ _3938_/Y _3926_/A _3939_/X _3933_/X VGND VGND VPWR VPWR _4957_/D sky130_fd_sc_hd__o211a_1
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3871_ _3597_/B _5038_/Q _3599_/B _5037_/Q VGND VGND VPWR VPWR _3871_/X sky130_fd_sc_hd__a211o_1
X_2822_ _4965_/Q _2787_/X _2788_/X VGND VGND VPWR VPWR _2830_/A sky130_fd_sc_hd__o21a_1
XFILLER_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2753_ _4965_/Q _2716_/X _2731_/X VGND VGND VPWR VPWR _2755_/C sky130_fd_sc_hd__o21a_1
X_2684_ _4942_/Q _2630_/B _2590_/C VGND VGND VPWR VPWR _2686_/C sky130_fd_sc_hd__o21a_1
X_4423_ _4410_/Y _4596_/A _4592_/A _4422_/X VGND VGND VPWR VPWR _4580_/A sky130_fd_sc_hd__o31a_1
X_4354_ _4326_/A _4848_/Q _4351_/X _4353_/Y VGND VGND VPWR VPWR _4354_/X sky130_fd_sc_hd__a22o_1
X_3305_ _3312_/A VGND VGND VPWR VPWR _3305_/X sky130_fd_sc_hd__buf_1
X_4285_ _4821_/Q _4285_/B VGND VGND VPWR VPWR _4285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3236_ _3340_/A _3008_/X _3235_/Y VGND VGND VPWR VPWR _3237_/B sky130_fd_sc_hd__o21ai_1
X_3167_ _3172_/A VGND VGND VPWR VPWR _3167_/X sky130_fd_sc_hd__buf_1
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3098_ _3098_/A VGND VGND VPWR VPWR _3308_/A sky130_fd_sc_hd__inv_2
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4070_ _4987_/Q VGND VGND VPWR VPWR _4070_/Y sky130_fd_sc_hd__inv_2
X_3021_ _5079_/Q _5116_/Q VGND VGND VPWR VPWR _3021_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4972_ _5018_/CLK _4972_/D VGND VGND VPWR VPWR _4972_/Q sky130_fd_sc_hd__dfxtp_1
X_3923_ _3923_/A _3923_/B VGND VGND VPWR VPWR _3924_/C sky130_fd_sc_hd__nand2_1
X_3854_ _3809_/A _3848_/Y _3809_/X _3852_/X _3853_/X VGND VGND VPWR VPWR _3854_/X
+ sky130_fd_sc_hd__o221a_1
X_2805_ _2721_/A _2774_/X _2775_/X VGND VGND VPWR VPWR _2807_/C sky130_fd_sc_hd__o21a_1
X_3785_ _3618_/B _5029_/Q _3618_/B _5029_/Q VGND VGND VPWR VPWR _3941_/A sky130_fd_sc_hd__a2bb2o_1
X_2736_ _2736_/A _2756_/B VGND VGND VPWR VPWR _2736_/X sky130_fd_sc_hd__or2_1
X_2667_ _4953_/Q VGND VGND VPWR VPWR _2746_/A sky130_fd_sc_hd__clkbuf_2
X_4406_ _4406_/A _4587_/B VGND VGND VPWR VPWR _4424_/C sky130_fd_sc_hd__nand2_1
X_2598_ _4967_/Q _4969_/Q _2615_/C VGND VGND VPWR VPWR _2611_/A sky130_fd_sc_hd__or3_4
XFILLER_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4337_ _4337_/A VGND VGND VPWR VPWR _4624_/B sky130_fd_sc_hd__clkbuf_2
X_4268_ _4268_/A VGND VGND VPWR VPWR _4268_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3219_ _3344_/A _2991_/X _3218_/Y VGND VGND VPWR VPWR _3220_/A sky130_fd_sc_hd__o21ai_1
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4199_ _4199_/A VGND VGND VPWR VPWR _4199_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3570_ _3478_/A _3478_/B _3568_/Y _3556_/A VGND VGND VPWR VPWR _5053_/D sky130_fd_sc_hd__a211oi_2
X_2521_ _4709_/B _2521_/B VGND VGND VPWR VPWR _2521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2452_ _4672_/A _2451_/B _2450_/X _2451_/Y VGND VGND VPWR VPWR _4815_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4122_ _4880_/Q _4053_/Y _3703_/B _4991_/Q VGND VGND VPWR VPWR _4123_/A sky130_fd_sc_hd__o22a_1
X_4053_ _4991_/Q VGND VGND VPWR VPWR _4053_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3004_ _3004_/A VGND VGND VPWR VPWR _3004_/X sky130_fd_sc_hd__clkbuf_2
Xinput3 dec_rate[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4955_ _5018_/CLK _4955_/D VGND VGND VPWR VPWR _4955_/Q sky130_fd_sc_hd__dfxtp_1
X_3906_ _3595_/B _5039_/Q _3905_/X VGND VGND VPWR VPWR _3907_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4886_ _5028_/CLK _4886_/D VGND VGND VPWR VPWR _4886_/Q sky130_fd_sc_hd__dfxtp_1
X_3837_ _5011_/Q VGND VGND VPWR VPWR _3837_/Y sky130_fd_sc_hd__inv_2
X_3768_ _3599_/B _5037_/Q _3599_/B _5037_/Q VGND VGND VPWR VPWR _3911_/A sky130_fd_sc_hd__a2bb2o_1
X_2719_ _2821_/A _2718_/X _2663_/X VGND VGND VPWR VPWR _2720_/D sky130_fd_sc_hd__o21a_1
X_3699_ _3703_/A _3699_/B VGND VGND VPWR VPWR _4993_/D sky130_fd_sc_hd__nor2_1
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4740_ _4740_/A _4740_/B _4740_/C _4740_/D VGND VGND VPWR VPWR _4740_/X sky130_fd_sc_hd__or4_4
X_4671_ _4458_/A _2972_/A _4814_/Q _5127_/Q VGND VGND VPWR VPWR _4672_/B sky130_fd_sc_hd__o22a_1
X_3622_ _3622_/A _3622_/B VGND VGND VPWR VPWR _5027_/D sky130_fd_sc_hd__nor2_1
X_3553_ _3556_/A VGND VGND VPWR VPWR _3559_/A sky130_fd_sc_hd__inv_2
X_3484_ _3484_/A _3484_/B VGND VGND VPWR VPWR _3562_/A sky130_fd_sc_hd__or2_1
X_2504_ _4706_/B _2512_/B _4743_/Y VGND VGND VPWR VPWR _2505_/B sky130_fd_sc_hd__o21ai_1
X_2435_ _4668_/B _2434_/B _2417_/X _2434_/Y VGND VGND VPWR VPWR _4819_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4105_ _3740_/B _4975_/Q _4864_/Q _4104_/Y VGND VGND VPWR VPWR _4105_/X sky130_fd_sc_hd__o22a_1
X_5085_ _3408_/X _5085_/D VGND VGND VPWR VPWR _5085_/Q sky130_fd_sc_hd__dfxtp_1
X_4036_ _4999_/Q VGND VGND VPWR VPWR _4036_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ _5018_/CLK _4938_/D VGND VGND VPWR VPWR _4938_/Q sky130_fd_sc_hd__dfxtp_1
X_4869_ _5018_/CLK _4869_/D VGND VGND VPWR VPWR _4869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2984_ _2984_/A _3207_/B VGND VGND VPWR VPWR _2985_/B sky130_fd_sc_hd__or2_1
X_4723_ _4793_/Q _5106_/Q _4721_/Y _4722_/Y VGND VGND VPWR VPWR _4724_/A sky130_fd_sc_hd__o22a_1
X_4654_ _4654_/A VGND VGND VPWR VPWR _4654_/Y sky130_fd_sc_hd__inv_2
X_3605_ _4923_/Q VGND VGND VPWR VPWR _3606_/B sky130_fd_sc_hd__inv_2
X_4585_ _4424_/A _4584_/Y _4391_/A _4584_/A _4575_/X VGND VGND VPWR VPWR _4870_/D
+ sky130_fd_sc_hd__o221a_1
X_3536_ _3516_/A _3516_/B _3517_/B VGND VGND VPWR VPWR _3536_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3467_ _4648_/A VGND VGND VPWR VPWR _3467_/X sky130_fd_sc_hd__buf_1
X_3398_ _5088_/Q _3397_/Y _3375_/X _3398_/C1 VGND VGND VPWR VPWR _5088_/D sky130_fd_sc_hd__o211a_1
X_2418_ _2416_/Y _4654_/A _2417_/X _2411_/X VGND VGND VPWR VPWR _4822_/D sky130_fd_sc_hd__o211a_1
X_5137_ _3172_/A _5137_/D VGND VGND VPWR VPWR _5137_/Q sky130_fd_sc_hd__dfxtp_1
X_5068_ _3455_/X _5068_/D VGND VGND VPWR VPWR _5068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4019_ _4019_/A VGND VGND VPWR VPWR _4019_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4370_ _4632_/B _4838_/Q _4369_/A _4838_/Q VGND VGND VPWR VPWR _4561_/A sky130_fd_sc_hd__a2bb2o_1
X_3321_ _3320_/X _3096_/B _5064_/Q _5101_/Q _3267_/X VGND VGND VPWR VPWR _5101_/D
+ sky130_fd_sc_hd__o221a_1
X_3252_ _3269_/A VGND VGND VPWR VPWR _3252_/X sky130_fd_sc_hd__buf_1
X_3183_ _3182_/A _3182_/B _3165_/X _3182_/Y VGND VGND VPWR VPWR _5132_/D sky130_fd_sc_hd__o211a_1
XFILLER_66_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2967_ _5128_/Q VGND VGND VPWR VPWR _2968_/A sky130_fd_sc_hd__inv_2
X_4706_ _4706_/A _4706_/B VGND VGND VPWR VPWR _4706_/X sky130_fd_sc_hd__or2_1
X_2898_ _5048_/Q VGND VGND VPWR VPWR _2903_/A sky130_fd_sc_hd__inv_2
X_4637_ _4638_/A _4637_/B VGND VGND VPWR VPWR _4834_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4568_ _4568_/A VGND VGND VPWR VPWR _4568_/Y sky130_fd_sc_hd__inv_2
X_4499_ _4499_/A VGND VGND VPWR VPWR _4499_/Y sky130_fd_sc_hd__inv_2
X_3519_ _2881_/A _3517_/X _3518_/X VGND VGND VPWR VPWR _3519_/X sky130_fd_sc_hd__a21bo_1
XFILLER_76_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3870_ _4925_/Q _3770_/Y _3869_/Y VGND VGND VPWR VPWR _3870_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2821_ _2821_/A _2821_/B VGND VGND VPWR VPWR _2821_/X sky130_fd_sc_hd__or2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2752_ _2752_/A _2752_/B _2752_/C _2752_/D VGND VGND VPWR VPWR _2755_/B sky130_fd_sc_hd__or4_4
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4422_ _4644_/B _4828_/Q _4408_/Y _4643_/B _4829_/Q VGND VGND VPWR VPWR _4422_/X
+ sky130_fd_sc_hd__o32a_1
X_2683_ _4939_/Q _2651_/X _2590_/B VGND VGND VPWR VPWR _2686_/B sky130_fd_sc_hd__o21a_1
X_4353_ _4327_/X _4328_/Y _4352_/Y VGND VGND VPWR VPWR _4353_/Y sky130_fd_sc_hd__o21ai_1
X_4284_ _4859_/Q VGND VGND VPWR VPWR _4285_/B sky130_fd_sc_hd__inv_2
X_3304_ _3072_/Y _3301_/Y _3080_/A _4578_/A _3303_/Y VGND VGND VPWR VPWR _5106_/D
+ sky130_fd_sc_hd__o311a_1
X_3235_ _3235_/A _3235_/B VGND VGND VPWR VPWR _3235_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3166_ _3163_/Y _2939_/A _3165_/X _3158_/X VGND VGND VPWR VPWR _5135_/D sky130_fd_sc_hd__o211a_1
X_3097_ _3090_/X _3091_/Y _3318_/B VGND VGND VPWR VPWR _3098_/A sky130_fd_sc_hd__o21ai_2
XFILLER_39_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3999_ _3994_/A _3994_/B _3978_/X _3995_/A VGND VGND VPWR VPWR _4941_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3020_ _3345_/A _2988_/Y _3344_/A _2991_/X _3019_/X VGND VGND VPWR VPWR _3020_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4971_ _5018_/CLK _4971_/D VGND VGND VPWR VPWR _4971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3922_ _3774_/A _3921_/Y _3772_/A _3921_/A _3902_/X VGND VGND VPWR VPWR _4962_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3853_ _3628_/B _5025_/Q _3799_/Y _3626_/B _5026_/Q VGND VGND VPWR VPWR _3853_/X
+ sky130_fd_sc_hd__o32a_1
X_2804_ _2680_/A _2791_/X _2772_/X VGND VGND VPWR VPWR _2807_/B sky130_fd_sc_hd__o21a_1
X_3784_ _3784_/A VGND VGND VPWR VPWR _3786_/A sky130_fd_sc_hd__inv_2
X_2735_ _2735_/A _2735_/B _2735_/C _2735_/D VGND VGND VPWR VPWR _2735_/X sky130_fd_sc_hd__or4_4
X_2666_ _2666_/A _2691_/B VGND VGND VPWR VPWR _2666_/X sky130_fd_sc_hd__or2_1
X_4405_ _4722_/A _4830_/Q _4398_/Y VGND VGND VPWR VPWR _4587_/B sky130_fd_sc_hd__a21oi_4
X_2597_ _4966_/Q _4965_/Q VGND VGND VPWR VPWR _2615_/C sky130_fd_sc_hd__or2_1
X_4336_ _4807_/Q VGND VGND VPWR VPWR _4337_/A sky130_fd_sc_hd__inv_2
X_4267_ _3736_/B _4976_/Q _4266_/X VGND VGND VPWR VPWR _4268_/A sky130_fd_sc_hd__o21ai_1
X_3218_ _3218_/A _3218_/B VGND VGND VPWR VPWR _3218_/Y sky130_fd_sc_hd__nand2_1
X_4198_ _3692_/B _4996_/Q _4197_/Y VGND VGND VPWR VPWR _4199_/A sky130_fd_sc_hd__o21ai_1
X_3149_ _2934_/Y _3158_/B _3163_/A _3148_/X VGND VGND VPWR VPWR _3150_/A sky130_fd_sc_hd__o31a_1
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2520_ _4741_/X _4715_/B _4745_/Y VGND VGND VPWR VPWR _2521_/B sky130_fd_sc_hd__o21ai_1
X_2451_ _4672_/A _2451_/B VGND VGND VPWR VPWR _2451_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4121_ _4075_/X _4084_/X _4250_/A _4120_/X VGND VGND VPWR VPWR _4219_/A sky130_fd_sc_hd__o31a_2
XFILLER_68_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4052_ _4052_/A _4208_/A VGND VGND VPWR VPWR _4127_/A sky130_fd_sc_hd__or2_1
X_3003_ _5120_/Q VGND VGND VPWR VPWR _3004_/A sky130_fd_sc_hd__inv_2
Xinput4 dec_rate[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4954_ _5018_/CLK _4954_/D VGND VGND VPWR VPWR _4954_/Q sky130_fd_sc_hd__dfxtp_1
X_3905_ _3909_/A _3905_/B VGND VGND VPWR VPWR _3905_/X sky130_fd_sc_hd__or2_1
X_4885_ _5028_/CLK _4885_/D VGND VGND VPWR VPWR _4885_/Q sky130_fd_sc_hd__dfxtp_1
X_3836_ _3654_/B _5013_/Q _3654_/B _5013_/Q VGND VGND VPWR VPWR _4004_/A sky130_fd_sc_hd__a2bb2o_1
X_3767_ _3597_/B _5038_/Q _3597_/B _5038_/Q VGND VGND VPWR VPWR _3916_/A sky130_fd_sc_hd__a2bb2o_1
X_2718_ _2783_/A VGND VGND VPWR VPWR _2718_/X sky130_fd_sc_hd__clkbuf_2
X_3698_ _4882_/Q VGND VGND VPWR VPWR _3699_/B sky130_fd_sc_hd__inv_2
X_2649_ _4943_/Q _2638_/X _2590_/A VGND VGND VPWR VPWR _2656_/A sky130_fd_sc_hd__o21a_1
X_4319_ _4319_/A _4517_/B VGND VGND VPWR VPWR _4320_/B sky130_fd_sc_hd__or2_1
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4670_ _4455_/A _2968_/A _4815_/Q _5128_/Q VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__o22a_1
X_3621_ _4916_/Q VGND VGND VPWR VPWR _3622_/B sky130_fd_sc_hd__inv_2
X_3552_ _2922_/A _2922_/B _3551_/X VGND VGND VPWR VPWR _3556_/A sky130_fd_sc_hd__o21ba_2
X_2503_ _2503_/A VGND VGND VPWR VPWR _2512_/B sky130_fd_sc_hd__inv_2
X_3483_ _3483_/A _3483_/B VGND VGND VPWR VPWR _3484_/B sky130_fd_sc_hd__nand2_1
X_2434_ _4668_/B _2434_/B VGND VGND VPWR VPWR _2434_/Y sky130_fd_sc_hd__nand2_1
X_4104_ _4975_/Q VGND VGND VPWR VPWR _4104_/Y sky130_fd_sc_hd__inv_2
X_5084_ _3410_/X _5084_/D VGND VGND VPWR VPWR _5084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4035_ _4184_/A _4179_/A VGND VGND VPWR VPWR _4041_/A sky130_fd_sc_hd__or2_1
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4937_ _5018_/CLK _4937_/D VGND VGND VPWR VPWR _4937_/Q sky130_fd_sc_hd__dfxtp_1
X_4868_ _5018_/CLK _4868_/D VGND VGND VPWR VPWR _4868_/Q sky130_fd_sc_hd__dfxtp_1
X_3819_ _5018_/Q VGND VGND VPWR VPWR _3820_/B sky130_fd_sc_hd__inv_2
X_4799_ _2519_/X _4799_/D VGND VGND VPWR VPWR _4799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2983_ _2983_/A VGND VGND VPWR VPWR _3207_/B sky130_fd_sc_hd__inv_2
X_4722_ _4722_/A _4722_/B VGND VGND VPWR VPWR _4722_/Y sky130_fd_sc_hd__nor2_4
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4653_ _4470_/A _2937_/A _4822_/Q _5135_/Q VGND VGND VPWR VPWR _4654_/A sky130_fd_sc_hd__o22a_1
X_3604_ _3611_/A _3604_/B VGND VGND VPWR VPWR _5035_/D sky130_fd_sc_hd__nor2_1
X_4584_ _4584_/A VGND VGND VPWR VPWR _4584_/Y sky130_fd_sc_hd__inv_2
X_3535_ _3525_/A _3525_/B _3525_/Y _3531_/X _3534_/X VGND VGND VPWR VPWR _3542_/A
+ sky130_fd_sc_hd__a2111o_1
X_3466_ _4647_/A _3466_/B _3466_/C VGND VGND VPWR VPWR _5066_/D sky130_fd_sc_hd__nor3_1
X_2417_ _3165_/A VGND VGND VPWR VPWR _2417_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3397_ _3397_/A VGND VGND VPWR VPWR _3397_/Y sky130_fd_sc_hd__inv_2
X_5136_ _3157_/X _5136_/D VGND VGND VPWR VPWR _5136_/Q sky130_fd_sc_hd__dfxtp_2
X_5067_ _3460_/X _5067_/D VGND VGND VPWR VPWR _5067_/Q sky130_fd_sc_hd__dfxtp_1
X_4018_ _4896_/Q _4017_/B _4017_/Y VGND VGND VPWR VPWR _4019_/A sky130_fd_sc_hd__a21oi_2
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3320_ _3324_/A VGND VGND VPWR VPWR _3320_/X sky130_fd_sc_hd__clkbuf_2
X_3251_ _3250_/Y _3123_/A _3223_/X _3242_/X VGND VGND VPWR VPWR _5117_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3182_ _3182_/A _3182_/B VGND VGND VPWR VPWR _3182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2966_ _5091_/Q VGND VGND VPWR VPWR _3349_/A sky130_fd_sc_hd__inv_1
X_2897_ _2897_/A VGND VGND VPWR VPWR _2897_/Y sky130_fd_sc_hd__inv_2
X_4705_ _4705_/A _4705_/B VGND VGND VPWR VPWR _4706_/B sky130_fd_sc_hd__or2_1
XFILLER_30_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4636_ _4638_/A _4636_/B VGND VGND VPWR VPWR _4835_/D sky130_fd_sc_hd__nor2_1
XFILLER_78_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4567_ _4635_/B _4836_/Q _4566_/Y VGND VGND VPWR VPWR _4568_/A sky130_fd_sc_hd__o21ai_1
X_4498_ _4613_/B _4854_/Q _4497_/X VGND VGND VPWR VPWR _4499_/A sky130_fd_sc_hd__o21ai_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3518_ _3518_/A _3518_/B VGND VGND VPWR VPWR _3518_/X sky130_fd_sc_hd__or2_1
X_3449_ _3329_/A _3449_/A2 _3431_/X _3446_/Y VGND VGND VPWR VPWR _5071_/D sky130_fd_sc_hd__a211oi_1
X_5119_ _3239_/X _5119_/D VGND VGND VPWR VPWR _5119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2820_ _2820_/A _2820_/B _2820_/C _2820_/D VGND VGND VPWR VPWR _2820_/X sky130_fd_sc_hd__or4_1
X_2751_ _2786_/A _2712_/X _2713_/X VGND VGND VPWR VPWR _2752_/D sky130_fd_sc_hd__o21a_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2682_ _2636_/B _2638_/X _2590_/A VGND VGND VPWR VPWR _2686_/A sky130_fd_sc_hd__o21a_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4421_ _4791_/Q VGND VGND VPWR VPWR _4643_/B sky130_fd_sc_hd__inv_2
X_4352_ _4622_/B _4847_/Q _4623_/B _4846_/Q VGND VGND VPWR VPWR _4352_/Y sky130_fd_sc_hd__o22ai_1
X_4283_ _4470_/A _4860_/Q _4470_/A _4860_/Q VGND VGND VPWR VPWR _4480_/B sky130_fd_sc_hd__a2bb2o_1
X_3303_ _3072_/Y _3301_/Y _3080_/A VGND VGND VPWR VPWR _3303_/Y sky130_fd_sc_hd__o21ai_1
X_3234_ _3250_/A _3125_/B _3013_/Y VGND VGND VPWR VPWR _3235_/B sky130_fd_sc_hd__o21ai_1
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3165_ _3165_/A VGND VGND VPWR VPWR _3165_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_66_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3096_ _3324_/A _3096_/B _3096_/C VGND VGND VPWR VPWR _3318_/B sky130_fd_sc_hd__or3_1
XFILLER_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3998_ _3825_/Y _3995_/Y _3831_/A _3996_/X _3997_/Y VGND VGND VPWR VPWR _4942_/D
+ sky130_fd_sc_hd__o311a_1
X_2949_ _5129_/Q VGND VGND VPWR VPWR _2949_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4619_ _4620_/A _4619_/B VGND VGND VPWR VPWR _4849_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4970_ _5018_/CLK _4970_/D VGND VGND VPWR VPWR _4970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3921_ _3921_/A VGND VGND VPWR VPWR _3921_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3852_ _3634_/B _5022_/Q _3818_/A _3850_/Y _3851_/X VGND VGND VPWR VPWR _3852_/X
+ sky130_fd_sc_hd__o221a_1
X_2803_ _4954_/Q _2770_/X _2758_/X VGND VGND VPWR VPWR _2807_/A sky130_fd_sc_hd__o21a_1
X_3783_ _3616_/B _5030_/Q _3616_/B _5030_/Q VGND VGND VPWR VPWR _3784_/A sky130_fd_sc_hd__o2bb2a_1
X_2734_ _2831_/A _2718_/X _2733_/X VGND VGND VPWR VPWR _2735_/D sky130_fd_sc_hd__o21a_1
X_2665_ _2665_/A _2665_/B _2665_/C _2665_/D VGND VGND VPWR VPWR _2665_/X sky130_fd_sc_hd__or4_1
X_2596_ _4957_/Q VGND VGND VPWR VPWR _2801_/A sky130_fd_sc_hd__clkbuf_2
X_4404_ _4721_/A _4831_/Q _4396_/Y VGND VGND VPWR VPWR _4406_/A sky130_fd_sc_hd__a21oi_4
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4335_ _4335_/A _4532_/A VGND VGND VPWR VPWR _4450_/C sky130_fd_sc_hd__or2_1
X_4266_ _4266_/A _4271_/A VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__or2_1
X_3217_ _3129_/C _3227_/B _3018_/Y VGND VGND VPWR VPWR _3218_/B sky130_fd_sc_hd__o21ai_1
X_4197_ _4197_/A _4197_/B VGND VGND VPWR VPWR _4197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3148_ _3356_/A _2937_/X _2932_/Y _3357_/A _3147_/Y VGND VGND VPWR VPWR _3148_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_54_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3079_ _3326_/A _4722_/B _3072_/Y VGND VGND VPWR VPWR _3300_/B sky130_fd_sc_hd__a21oi_4
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2450_ _3165_/A VGND VGND VPWR VPWR _2450_/X sky130_fd_sc_hd__buf_2
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4120_ _4075_/A _4114_/Y _4075_/X _4118_/X _4119_/X VGND VGND VPWR VPWR _4120_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4051_ _3701_/B _4992_/Q _3701_/B _4992_/Q VGND VGND VPWR VPWR _4208_/A sky130_fd_sc_hd__a2bb2o_1
Xinput5 dec_rate[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_2
X_3002_ _5083_/Q VGND VGND VPWR VPWR _3341_/A sky130_fd_sc_hd__inv_1
XFILLER_76_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4953_ _5018_/CLK _4953_/D VGND VGND VPWR VPWR _4953_/Q sky130_fd_sc_hd__dfxtp_1
X_3904_ _3899_/A _3899_/B _3462_/X _3899_/Y VGND VGND VPWR VPWR _4967_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4884_ _5028_/CLK _4884_/D VGND VGND VPWR VPWR _4884_/Q sky130_fd_sc_hd__dfxtp_1
X_3835_ _3835_/A VGND VGND VPWR VPWR _3835_/Y sky130_fd_sc_hd__inv_2
X_3766_ _3766_/A _3766_/B VGND VGND VPWR VPWR _3766_/X sky130_fd_sc_hd__or2_1
X_2717_ _4962_/Q _2716_/X _2659_/X VGND VGND VPWR VPWR _2720_/C sky130_fd_sc_hd__o21a_1
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3697_ _3703_/A _3697_/B VGND VGND VPWR VPWR _4994_/D sky130_fd_sc_hd__nor2_1
X_2648_ _2736_/A _2645_/X _2647_/X VGND VGND VPWR VPWR _2665_/A sky130_fd_sc_hd__o21a_1
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2579_ _2758_/A VGND VGND VPWR VPWR _2590_/A sky130_fd_sc_hd__buf_1
X_4318_ _4618_/B _4850_/Q _4317_/A _4850_/Q VGND VGND VPWR VPWR _4517_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4249_ _4083_/A _4248_/Y _4081_/A _4248_/A _4229_/X VGND VGND VPWR VPWR _4909_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3620_ _3622_/A _3620_/B VGND VGND VPWR VPWR _5028_/D sky130_fd_sc_hd__nor2_1
X_3551_ _3551_/A _3551_/B _3550_/X VGND VGND VPWR VPWR _3551_/X sky130_fd_sc_hd__or3b_2
X_2502_ _4741_/X _4715_/X _4747_/X VGND VGND VPWR VPWR _2503_/A sky130_fd_sc_hd__o21ai_1
X_3482_ _3482_/A VGND VGND VPWR VPWR _3483_/B sky130_fd_sc_hd__inv_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2433_ _4611_/B _2960_/X _2432_/Y VGND VGND VPWR VPWR _2434_/B sky130_fd_sc_hd__o21ai_1
X_4103_ _4974_/Q VGND VGND VPWR VPWR _4103_/Y sky130_fd_sc_hd__inv_2
X_5083_ _3413_/X _5083_/D VGND VGND VPWR VPWR _5083_/Q sky130_fd_sc_hd__dfxtp_1
X_4034_ _3683_/B _5000_/Q _3683_/B _5000_/Q VGND VGND VPWR VPWR _4179_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4936_ _5047_/CLK _4936_/D VGND VGND VPWR VPWR _4936_/Q sky130_fd_sc_hd__dfxtp_1
X_4867_ _5018_/CLK _4867_/D VGND VGND VPWR VPWR _4867_/Q sky130_fd_sc_hd__dfxtp_1
X_3818_ _3818_/A _3818_/B VGND VGND VPWR VPWR _3818_/X sky130_fd_sc_hd__or2_1
X_4798_ _2526_/X _4798_/D VGND VGND VPWR VPWR _4798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3749_ _3582_/B _5045_/Q _3582_/B _5045_/Q VGND VGND VPWR VPWR _3887_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2982_ _3346_/A _2981_/Y _5088_/Q _5125_/Q VGND VGND VPWR VPWR _2983_/A sky130_fd_sc_hd__o22a_1
XFILLER_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4721_ _4721_/A _4721_/B VGND VGND VPWR VPWR _4721_/Y sky130_fd_sc_hd__nor2_2
X_4652_ _4652_/A VGND VGND VPWR VPWR _4652_/Y sky130_fd_sc_hd__inv_2
X_3603_ _4924_/Q VGND VGND VPWR VPWR _3604_/B sky130_fd_sc_hd__inv_2
X_4583_ _4640_/B _4832_/Q _4582_/Y VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__o21ai_1
X_3534_ _2910_/X _3533_/X _2910_/X _3533_/X VGND VGND VPWR VPWR _3534_/X sky130_fd_sc_hd__a2bb2o_1
X_3465_ _3320_/X _3465_/A2 _3090_/X _3324_/D VGND VGND VPWR VPWR _3466_/C sky130_fd_sc_hd__o31a_1
X_2416_ _2416_/A VGND VGND VPWR VPWR _2416_/Y sky130_fd_sc_hd__inv_2
X_3396_ _3396_/A VGND VGND VPWR VPWR _3396_/X sky130_fd_sc_hd__buf_1
X_5135_ _3162_/X _5135_/D VGND VGND VPWR VPWR _5135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5066_ _3464_/X _5066_/D VGND VGND VPWR VPWR _5066_/Q sky130_fd_sc_hd__dfxtp_1
X_4017_ _4896_/Q _4017_/B VGND VGND VPWR VPWR _4017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4919_ _5047_/CLK _4919_/D VGND VGND VPWR VPWR _4919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3250_ _3250_/A VGND VGND VPWR VPWR _3250_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3181_ _3352_/A _2960_/X _3180_/Y VGND VGND VPWR VPWR _3182_/B sky130_fd_sc_hd__o21ai_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4704_ _4704_/A VGND VGND VPWR VPWR _4705_/B sky130_fd_sc_hd__inv_2
X_2965_ _2965_/A _2965_/B VGND VGND VPWR VPWR _2965_/X sky130_fd_sc_hd__or2_1
X_2896_ _3523_/A _2845_/B _2846_/B VGND VGND VPWR VPWR _2897_/A sky130_fd_sc_hd__a21bo_1
X_4635_ _4638_/A _4635_/B VGND VGND VPWR VPWR _4836_/D sky130_fd_sc_hd__nor2_1
X_4566_ _4566_/A _4566_/B VGND VGND VPWR VPWR _4566_/Y sky130_fd_sc_hd__nand2_1
X_3517_ _3517_/A _3517_/B VGND VGND VPWR VPWR _3517_/X sky130_fd_sc_hd__or2_2
X_4497_ _4503_/A _4497_/B VGND VGND VPWR VPWR _4497_/X sky130_fd_sc_hd__or2_1
X_3448_ _3455_/A VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__buf_1
X_3379_ _3382_/A VGND VGND VPWR VPWR _3379_/X sky130_fd_sc_hd__buf_1
XFILLER_69_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5118_ _3241_/X _5118_/D VGND VGND VPWR VPWR _5118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5049_ _5063_/CLK _5049_/D VGND VGND VPWR VPWR _5049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ _2666_/A _2709_/X _2710_/X VGND VGND VPWR VPWR _2752_/C sky130_fd_sc_hd__o21a_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2681_ _2756_/A _2645_/X _2647_/X VGND VGND VPWR VPWR _2690_/A sky130_fd_sc_hd__o21a_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4420_ _4420_/A VGND VGND VPWR VPWR _4644_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4351_ _4450_/C _4351_/B VGND VGND VPWR VPWR _4351_/X sky130_fd_sc_hd__or2_1
X_3302_ _4153_/A VGND VGND VPWR VPWR _4578_/A sky130_fd_sc_hd__clkbuf_4
X_4282_ _4822_/Q VGND VGND VPWR VPWR _4470_/A sky130_fd_sc_hd__inv_2
X_3233_ _3241_/A VGND VGND VPWR VPWR _3233_/X sky130_fd_sc_hd__buf_1
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3164_ _4176_/A VGND VGND VPWR VPWR _3165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3095_ _5065_/Q _5102_/Q _3090_/X _3091_/Y VGND VGND VPWR VPWR _3096_/C sky130_fd_sc_hd__a22o_1
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3997_ _3825_/Y _3995_/Y _3831_/A VGND VGND VPWR VPWR _3997_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2948_ _5092_/Q VGND VGND VPWR VPWR _3350_/A sky130_fd_sc_hd__clkinv_1
X_4618_ _4620_/A _4618_/B VGND VGND VPWR VPWR _4850_/D sky130_fd_sc_hd__nor2_1
X_2879_ _2879_/A VGND VGND VPWR VPWR _2879_/Y sky130_fd_sc_hd__inv_2
X_4549_ _4577_/A _4387_/X _4433_/X VGND VGND VPWR VPWR _4550_/A sky130_fd_sc_hd__o21ai_1
XFILLER_38_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3920_ _3604_/B _5035_/Q _3924_/B VGND VGND VPWR VPWR _3921_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3851_ _3634_/B _5022_/Q _3637_/B _5021_/Q VGND VGND VPWR VPWR _3851_/X sky130_fd_sc_hd__a211o_1
X_2802_ _4963_/Q _2787_/X _2788_/X VGND VGND VPWR VPWR _2810_/A sky130_fd_sc_hd__o21a_1
X_3782_ _3782_/A _3938_/A VGND VGND VPWR VPWR _3865_/C sky130_fd_sc_hd__or2_1
X_2733_ _2798_/A VGND VGND VPWR VPWR _2733_/X sky130_fd_sc_hd__buf_1
X_2664_ _2768_/A _2613_/B _2663_/X VGND VGND VPWR VPWR _2665_/D sky130_fd_sc_hd__o21a_1
X_4403_ _4640_/B _4832_/Q _4389_/Y _4638_/B _4833_/Q VGND VGND VPWR VPWR _4403_/X
+ sky130_fd_sc_hd__o32a_1
X_2595_ _2590_/X _2646_/A _2658_/A _2662_/A VGND VGND VPWR VPWR _4770_/S sky130_fd_sc_hd__and4b_4
X_4334_ _4623_/B _4846_/Q _4333_/A _4846_/Q VGND VGND VPWR VPWR _4532_/A sky130_fd_sc_hd__a2bb2o_1
X_4265_ _4260_/A _4260_/B _4264_/X _4261_/A VGND VGND VPWR VPWR _4904_/D sky130_fd_sc_hd__o211a_1
X_3216_ _3216_/A VGND VGND VPWR VPWR _3227_/B sky130_fd_sc_hd__inv_2
X_4196_ _4131_/C _4202_/B _4061_/Y VGND VGND VPWR VPWR _4197_/B sky130_fd_sc_hd__o21ai_1
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3147_ _5136_/Q VGND VGND VPWR VPWR _3147_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3078_ _3327_/A _4721_/B _3069_/Y VGND VGND VPWR VPWR _3080_/A sky130_fd_sc_hd__a21oi_4
XFILLER_35_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4050_ _4050_/A VGND VGND VPWR VPWR _4052_/A sky130_fd_sc_hd__inv_2
XFILLER_49_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3001_ _3001_/A _3227_/A VGND VGND VPWR VPWR _3129_/C sky130_fd_sc_hd__or2_1
Xinput6 dec_rate[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__buf_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4952_ _5018_/CLK _4952_/D VGND VGND VPWR VPWR _4952_/Q sky130_fd_sc_hd__dfxtp_1
X_3903_ _3765_/B _3901_/Y _3764_/A _3901_/A _3902_/X VGND VGND VPWR VPWR _4968_/D
+ sky130_fd_sc_hd__o221a_1
X_4883_ _5028_/CLK _4883_/D VGND VGND VPWR VPWR _4883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3834_ _4903_/Q _3833_/B _3833_/Y VGND VGND VPWR VPWR _3835_/A sky130_fd_sc_hd__a21oi_2
X_3765_ _3895_/A _3765_/B VGND VGND VPWR VPWR _3766_/B sky130_fd_sc_hd__or2_1
X_2716_ _2781_/A VGND VGND VPWR VPWR _2716_/X sky130_fd_sc_hd__clkbuf_2
X_3696_ _4883_/Q VGND VGND VPWR VPWR _3697_/B sky130_fd_sc_hd__inv_2
X_2647_ _2788_/A VGND VGND VPWR VPWR _2647_/X sky130_fd_sc_hd__buf_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2578_ _2881_/Y _2580_/B _3517_/X VGND VGND VPWR VPWR _2758_/A sky130_fd_sc_hd__nor3_4
X_4317_ _4317_/A VGND VGND VPWR VPWR _4618_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4248_ _4248_/A VGND VGND VPWR VPWR _4248_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4179_ _4179_/A VGND VGND VPWR VPWR _4181_/A sky130_fd_sc_hd__inv_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3550_ _5061_/Q _3546_/Y _3485_/A _3514_/X _3549_/Y VGND VGND VPWR VPWR _3550_/X
+ sky130_fd_sc_hd__o221a_1
X_2501_ _2519_/A VGND VGND VPWR VPWR _2501_/X sky130_fd_sc_hd__buf_1
X_3481_ _3481_/A _3481_/B VGND VGND VPWR VPWR _3482_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2432_ _4668_/A _2432_/B VGND VGND VPWR VPWR _2432_/Y sky130_fd_sc_hd__nand2_1
X_5082_ _3416_/X _5082_/D VGND VGND VPWR VPWR _5082_/Q sky130_fd_sc_hd__dfxtp_1
X_4102_ _3736_/B _4976_/Q _3736_/B _4976_/Q VGND VGND VPWR VPWR _4271_/A sky130_fd_sc_hd__a2bb2o_1
X_4033_ _3679_/B _5001_/Q _3679_/B _5001_/Q VGND VGND VPWR VPWR _4184_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4935_ _5047_/CLK _4935_/D VGND VGND VPWR VPWR _4935_/Q sky130_fd_sc_hd__dfxtp_1
X_4866_ _5018_/CLK _4866_/D VGND VGND VPWR VPWR _4866_/Q sky130_fd_sc_hd__dfxtp_1
X_4797_ _2528_/X _4797_/D VGND VGND VPWR VPWR _4797_/Q sky130_fd_sc_hd__dfxtp_1
X_3817_ _3817_/A _3984_/B VGND VGND VPWR VPWR _3818_/B sky130_fd_sc_hd__or2_1
X_3748_ _3748_/A VGND VGND VPWR VPWR _3748_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3679_ _3679_/A _3679_/B VGND VGND VPWR VPWR _5001_/D sky130_fd_sc_hd__nor2_1
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2981_ _5125_/Q VGND VGND VPWR VPWR _2981_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4720_ _4720_/A VGND VGND VPWR VPWR _4740_/B sky130_fd_sc_hd__inv_2
X_4651_ _4823_/Q _5136_/Q _4650_/Y VGND VGND VPWR VPWR _4652_/A sky130_fd_sc_hd__a21oi_2
X_3602_ _3611_/A _3602_/B VGND VGND VPWR VPWR _5036_/D sky130_fd_sc_hd__nor2_1
X_4582_ _4582_/A _4582_/B VGND VGND VPWR VPWR _4582_/Y sky130_fd_sc_hd__nand2_1
X_3533_ _3532_/Y _3523_/Y _3516_/B VGND VGND VPWR VPWR _3533_/X sky130_fd_sc_hd__o21a_1
X_3464_ _4648_/A VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__buf_1
X_2415_ _2428_/A VGND VGND VPWR VPWR _2415_/X sky130_fd_sc_hd__buf_1
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3395_ _3347_/A _3395_/A2 _3371_/X _3392_/Y VGND VGND VPWR VPWR _5089_/D sky130_fd_sc_hd__a211oi_1
X_5134_ _3167_/X _5134_/D VGND VGND VPWR VPWR _5134_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5065_ _3467_/X _5065_/D VGND VGND VPWR VPWR _5065_/Q sky130_fd_sc_hd__dfxtp_1
X_4016_ _5007_/Q VGND VGND VPWR VPWR _4017_/B sky130_fd_sc_hd__inv_2
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4918_ _5028_/CLK _4918_/D VGND VGND VPWR VPWR _4918_/Q sky130_fd_sc_hd__dfxtp_1
X_4849_ _5028_/CLK _4849_/D VGND VGND VPWR VPWR _4849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3180_ _3180_/A _3180_/B VGND VGND VPWR VPWR _3180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2964_ _3180_/A _3182_/A VGND VGND VPWR VPWR _2965_/B sky130_fd_sc_hd__nand2_1
X_4703_ _4369_/A _3034_/Y _4800_/Q _5113_/Q VGND VGND VPWR VPWR _4704_/A sky130_fd_sc_hd__o22a_1
X_2895_ _5050_/Q VGND VGND VPWR VPWR _2895_/Y sky130_fd_sc_hd__inv_2
X_4634_ _4638_/A _4634_/B VGND VGND VPWR VPWR _4837_/D sky130_fd_sc_hd__nor2_1
X_4565_ _4577_/A _4387_/B _4430_/Y VGND VGND VPWR VPWR _4566_/B sky130_fd_sc_hd__o21ai_1
X_3516_ _3516_/A _3516_/B VGND VGND VPWR VPWR _3517_/B sky130_fd_sc_hd__or2_1
X_4496_ _4492_/A _4492_/B _4264_/X _4492_/Y VGND VGND VPWR VPWR _4893_/D sky130_fd_sc_hd__o211a_1
X_3447_ _5072_/Q _3446_/Y _3435_/X _3447_/C1 VGND VGND VPWR VPWR _5072_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3378_ _3353_/A _3378_/A2 _3371_/X _3374_/Y VGND VGND VPWR VPWR _5095_/D sky130_fd_sc_hd__a211oi_1
XFILLER_57_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5117_ _3249_/X _5117_/D VGND VGND VPWR VPWR _5117_/Q sky130_fd_sc_hd__dfxtp_1
X_5048_ _5063_/CLK _5048_/D VGND VGND VPWR VPWR _5048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _2680_/A _2691_/B VGND VGND VPWR VPWR _2680_/X sky130_fd_sc_hd__or2_1
X_4350_ _4624_/B _4845_/Q _4446_/A _4347_/Y _4349_/X VGND VGND VPWR VPWR _4351_/B
+ sky130_fd_sc_hd__o221a_1
X_3301_ _3301_/A VGND VGND VPWR VPWR _3301_/Y sky130_fd_sc_hd__inv_2
X_4281_ _4281_/A VGND VGND VPWR VPWR _4281_/Y sky130_fd_sc_hd__inv_2
X_3232_ _3000_/A _3216_/A _3223_/X _3227_/X VGND VGND VPWR VPWR _5121_/D sky130_fd_sc_hd__o211a_1
X_3163_ _3163_/A VGND VGND VPWR VPWR _3163_/Y sky130_fd_sc_hd__inv_2
X_3094_ _4735_/B VGND VGND VPWR VPWR _3096_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3996_ _4153_/A VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__buf_2
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2947_ _2947_/A VGND VGND VPWR VPWR _3168_/B sky130_fd_sc_hd__inv_2
X_4617_ _4620_/A _4617_/B VGND VGND VPWR VPWR _4851_/D sky130_fd_sc_hd__nor2_1
X_2878_ input4/X _3507_/B _3508_/B VGND VGND VPWR VPWR _2879_/A sky130_fd_sc_hd__a21bo_1
X_4548_ _4548_/A VGND VGND VPWR VPWR _4552_/A sky130_fd_sc_hd__inv_2
X_4479_ _4281_/Y _4478_/Y _4281_/A _4478_/A _4269_/X VGND VGND VPWR VPWR _4898_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3850_ _4909_/Q _3813_/Y _3849_/Y VGND VGND VPWR VPWR _3850_/Y sky130_fd_sc_hd__o21ai_1
X_2801_ _2801_/A _2821_/B VGND VGND VPWR VPWR _2801_/X sky130_fd_sc_hd__or2_1
X_3781_ _3614_/B _5031_/Q _3614_/B _5031_/Q VGND VGND VPWR VPWR _3938_/A sky130_fd_sc_hd__a2bb2o_1
X_2732_ _4963_/Q _2716_/X _2731_/X VGND VGND VPWR VPWR _2735_/C sky130_fd_sc_hd__o21a_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2663_ _2798_/A VGND VGND VPWR VPWR _2663_/X sky130_fd_sc_hd__buf_1
X_4402_ _4795_/Q VGND VGND VPWR VPWR _4638_/B sky130_fd_sc_hd__inv_2
X_2594_ _2864_/Y _3513_/A _2858_/A VGND VGND VPWR VPWR _2662_/A sky130_fd_sc_hd__or3_4
X_4333_ _4333_/A VGND VGND VPWR VPWR _4623_/B sky130_fd_sc_hd__buf_1
XFILLER_59_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4264_ _4562_/A VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__clkbuf_4
X_3215_ _3250_/A _3129_/A _3016_/B VGND VGND VPWR VPWR _3216_/A sky130_fd_sc_hd__o21ai_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4195_ _4195_/A VGND VGND VPWR VPWR _4202_/B sky130_fd_sc_hd__inv_2
X_3146_ _5099_/Q VGND VGND VPWR VPWR _3357_/A sky130_fd_sc_hd__inv_2
X_3077_ _3328_/A _3064_/X _3059_/Y _3329_/A _3076_/Y VGND VGND VPWR VPWR _3077_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3979_ _3971_/A _3971_/B _3978_/X _3971_/Y VGND VGND VPWR VPWR _4947_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3000_ _3000_/A VGND VGND VPWR VPWR _3227_/A sky130_fd_sc_hd__inv_2
Xinput7 dec_rate[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4951_ _5018_/CLK _4951_/D VGND VGND VPWR VPWR _4951_/Q sky130_fd_sc_hd__dfxtp_1
X_4882_ _5028_/CLK _4882_/D VGND VGND VPWR VPWR _4882_/Q sky130_fd_sc_hd__dfxtp_1
X_3902_ _3936_/A VGND VGND VPWR VPWR _3902_/X sky130_fd_sc_hd__clkbuf_2
X_3833_ _4903_/Q _3833_/B VGND VGND VPWR VPWR _3833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3764_ _3764_/A VGND VGND VPWR VPWR _3765_/B sky130_fd_sc_hd__inv_2
X_2715_ _2715_/A _2715_/B _2715_/C _2715_/D VGND VGND VPWR VPWR _2720_/B sky130_fd_sc_hd__or4_4
X_3695_ _3703_/A _3695_/B VGND VGND VPWR VPWR _4995_/D sky130_fd_sc_hd__nor2_1
X_2646_ _2646_/A VGND VGND VPWR VPWR _2788_/A sky130_fd_sc_hd__inv_2
X_2577_ _2850_/A _3501_/A _2587_/D VGND VGND VPWR VPWR _2580_/B sky130_fd_sc_hd__or3_4
XFILLER_59_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4316_ _4812_/Q VGND VGND VPWR VPWR _4317_/A sky130_fd_sc_hd__inv_2
X_4247_ _3723_/B _4982_/Q _4251_/B VGND VGND VPWR VPWR _4248_/A sky130_fd_sc_hd__o21ai_1
X_4178_ _4175_/Y _4164_/A _4177_/X _4171_/X VGND VGND VPWR VPWR _4928_/D sky130_fd_sc_hd__o211a_1
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3129_ _3129_/A _3129_/B _3129_/C _3218_/A VGND VGND VPWR VPWR _3129_/X sky130_fd_sc_hd__or4b_4
XFILLER_55_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3480_ _3480_/A _3480_/B VGND VGND VPWR VPWR _3481_/B sky130_fd_sc_hd__nor2_2
X_2500_ _3384_/A VGND VGND VPWR VPWR _2519_/A sky130_fd_sc_hd__buf_1
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2431_ _4669_/A _2440_/B _2394_/Y VGND VGND VPWR VPWR _2432_/B sky130_fd_sc_hd__o21ai_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5081_ _3419_/X _5081_/D VGND VGND VPWR VPWR _5081_/Q sky130_fd_sc_hd__dfxtp_1
X_4101_ _4101_/A VGND VGND VPWR VPWR _4101_/Y sky130_fd_sc_hd__inv_2
X_4032_ _4032_/A _4032_/B VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__or2_1
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4934_ _5047_/CLK _4934_/D VGND VGND VPWR VPWR _4934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4865_ _5018_/CLK _4865_/D VGND VGND VPWR VPWR _4865_/Q sky130_fd_sc_hd__dfxtp_1
X_4796_ _2533_/X _4796_/D VGND VGND VPWR VPWR _4796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3816_ _3641_/B _5019_/Q _3641_/B _5019_/Q VGND VGND VPWR VPWR _3984_/B sky130_fd_sc_hd__a2bb2o_1
X_3747_ _4935_/Q _3746_/B _3746_/Y VGND VGND VPWR VPWR _3748_/A sky130_fd_sc_hd__a21oi_2
X_3678_ _4890_/Q VGND VGND VPWR VPWR _3679_/B sky130_fd_sc_hd__inv_2
X_2629_ _2774_/A VGND VGND VPWR VPWR _2630_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2980_ _5088_/Q VGND VGND VPWR VPWR _3346_/A sky130_fd_sc_hd__clkinv_1
XFILLER_42_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4650_ _4823_/Q _5136_/Q VGND VGND VPWR VPWR _4650_/Y sky130_fd_sc_hd__nor2_1
X_3601_ _4925_/Q VGND VGND VPWR VPWR _3602_/B sky130_fd_sc_hd__inv_2
Xinput10 dec_rate[3] VGND VGND VPWR VPWR _3523_/A sky130_fd_sc_hd__clkbuf_2
X_4581_ _4406_/A _4587_/B _4587_/A _4400_/A VGND VGND VPWR VPWR _4582_/B sky130_fd_sc_hd__a31o_1
X_3532_ _3532_/A VGND VGND VPWR VPWR _3532_/Y sky130_fd_sc_hd__inv_2
X_3463_ _5067_/Q _3466_/B _3462_/X _3463_/C1 VGND VGND VPWR VPWR _5067_/D sky130_fd_sc_hd__o211a_1
X_2414_ _4652_/Y _2413_/Y _4652_/A _2413_/A _4575_/X VGND VGND VPWR VPWR _4823_/D
+ sky130_fd_sc_hd__o221a_1
X_3394_ _3396_/A VGND VGND VPWR VPWR _3394_/X sky130_fd_sc_hd__buf_1
X_5133_ _3172_/X _5133_/D VGND VGND VPWR VPWR _5133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5064_ _3470_/X _5064_/D VGND VGND VPWR VPWR _5064_/Q sky130_fd_sc_hd__dfxtp_1
X_4015_ _3664_/B _5008_/Q _3664_/B _5008_/Q VGND VGND VPWR VPWR _4154_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4917_ _5028_/CLK _4917_/D VGND VGND VPWR VPWR _4917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4848_ _5028_/CLK _4848_/D VGND VGND VPWR VPWR _4848_/Q sky130_fd_sc_hd__dfxtp_1
X_4779_ _5139_/Q _4779_/D VGND VGND VPWR VPWR _4779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2963_ _5095_/Q _5132_/Q _2962_/Y VGND VGND VPWR VPWR _3182_/A sky130_fd_sc_hd__a21oi_2
X_4702_ _4702_/A VGND VGND VPWR VPWR _4705_/A sky130_fd_sc_hd__inv_2
X_2894_ _2894_/A VGND VGND VPWR VPWR _2894_/Y sky130_fd_sc_hd__inv_2
X_4633_ _4639_/A VGND VGND VPWR VPWR _4638_/A sky130_fd_sc_hd__clkbuf_2
X_4564_ _4564_/A VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__inv_2
X_3515_ _3518_/A _3515_/B VGND VGND VPWR VPWR _3516_/B sky130_fd_sc_hd__or2_2
X_4495_ _4304_/B _4494_/Y _4303_/A _4494_/A _4269_/X VGND VGND VPWR VPWR _4894_/D
+ sky130_fd_sc_hd__o221a_1
X_3446_ _3446_/A VGND VGND VPWR VPWR _3446_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3377_ _3382_/A VGND VGND VPWR VPWR _3377_/X sky130_fd_sc_hd__buf_1
X_5116_ _3252_/X _5116_/D VGND VGND VPWR VPWR _5116_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5047_ _5047_/CLK _5047_/D VGND VGND VPWR VPWR _5047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3300_ _3300_/A _3300_/B VGND VGND VPWR VPWR _3301_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4280_ _4823_/Q _4279_/B _4279_/Y VGND VGND VPWR VPWR _4281_/A sky130_fd_sc_hd__a21oi_2
X_3231_ _3241_/A VGND VGND VPWR VPWR _3231_/X sky130_fd_sc_hd__buf_1
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3162_ _3172_/A VGND VGND VPWR VPWR _3162_/X sky130_fd_sc_hd__buf_1
XFILLER_66_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3093_ _5101_/Q VGND VGND VPWR VPWR _4735_/B sky130_fd_sc_hd__inv_2
XFILLER_62_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_mclk1 clkbuf_0_mclk1/X VGND VGND VPWR VPWR _5063_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3995_ _3995_/A VGND VGND VPWR VPWR _3995_/Y sky130_fd_sc_hd__inv_2
X_2946_ _3354_/A _2945_/X _5096_/Q _5133_/Q VGND VGND VPWR VPWR _2947_/A sky130_fd_sc_hd__o22a_1
X_2877_ _5059_/Q VGND VGND VPWR VPWR _3485_/A sky130_fd_sc_hd__inv_2
X_4616_ _4620_/A _4616_/B VGND VGND VPWR VPWR _4852_/D sky130_fd_sc_hd__nor2_1
X_4547_ _4546_/Y _4444_/A _4526_/X _4542_/X VGND VGND VPWR VPWR _4879_/D sky130_fd_sc_hd__o211a_1
X_4478_ _4478_/A VGND VGND VPWR VPWR _4478_/Y sky130_fd_sc_hd__inv_2
X_3429_ _3444_/A VGND VGND VPWR VPWR _3442_/A sky130_fd_sc_hd__buf_1
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2800_ _2800_/A _2800_/B _2800_/C _2800_/D VGND VGND VPWR VPWR _2800_/X sky130_fd_sc_hd__or4_1
X_3780_ _3780_/A VGND VGND VPWR VPWR _3782_/A sky130_fd_sc_hd__inv_2
X_2731_ _2796_/A VGND VGND VPWR VPWR _2731_/X sky130_fd_sc_hd__buf_1
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2662_ _2662_/A VGND VGND VPWR VPWR _2798_/A sky130_fd_sc_hd__inv_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4401_ _4401_/A VGND VGND VPWR VPWR _4640_/B sky130_fd_sc_hd__clkbuf_2
X_2593_ _3498_/A _3507_/B _2593_/C VGND VGND VPWR VPWR _2658_/A sky130_fd_sc_hd__or3_4
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4332_ _4808_/Q VGND VGND VPWR VPWR _4333_/A sky130_fd_sc_hd__inv_2
X_4263_ _4091_/Y _4261_/Y _4097_/A _3996_/X _4262_/Y VGND VGND VPWR VPWR _4905_/D
+ sky130_fd_sc_hd__o311a_1
X_3214_ _3222_/A VGND VGND VPWR VPWR _3214_/X sky130_fd_sc_hd__buf_1
XFILLER_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4194_ _4219_/A _4131_/A _4059_/B VGND VGND VPWR VPWR _4195_/A sky130_fd_sc_hd__o21ai_1
X_3145_ _2942_/Y _3168_/B _3173_/A _3144_/X VGND VGND VPWR VPWR _3163_/A sky130_fd_sc_hd__o31a_1
X_3076_ _5108_/Q VGND VGND VPWR VPWR _3076_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3978_ _3978_/A VGND VGND VPWR VPWR _3978_/X sky130_fd_sc_hd__buf_2
X_2929_ _5100_/Q VGND VGND VPWR VPWR _2929_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_40_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 dec_rate[1] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4950_ _5018_/CLK _4950_/D VGND VGND VPWR VPWR _4950_/Q sky130_fd_sc_hd__dfxtp_1
X_3901_ _3901_/A VGND VGND VPWR VPWR _3901_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4881_ _5028_/CLK _4881_/D VGND VGND VPWR VPWR _4881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3832_ _5014_/Q VGND VGND VPWR VPWR _3833_/B sky130_fd_sc_hd__inv_2
X_3763_ _4931_/Q _3762_/B _3762_/Y VGND VGND VPWR VPWR _3764_/A sky130_fd_sc_hd__a21oi_2
X_2714_ _2746_/A _2712_/X _2713_/X VGND VGND VPWR VPWR _2715_/D sky130_fd_sc_hd__o21a_1
X_3694_ _4884_/Q VGND VGND VPWR VPWR _3695_/B sky130_fd_sc_hd__inv_2
X_2645_ _2787_/A VGND VGND VPWR VPWR _2645_/X sky130_fd_sc_hd__buf_1
X_4315_ _4315_/A VGND VGND VPWR VPWR _4319_/A sky130_fd_sc_hd__inv_2
X_2576_ _2866_/A input3/X _2858_/A VGND VGND VPWR VPWR _2587_/D sky130_fd_sc_hd__or3_1
XFILLER_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4246_ _4250_/A _4250_/B VGND VGND VPWR VPWR _4251_/B sky130_fd_sc_hd__or2_1
X_4177_ _4562_/A VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__clkbuf_2
X_3128_ _5086_/Q _5123_/Q _3344_/A _2991_/A VGND VGND VPWR VPWR _3218_/A sky130_fd_sc_hd__o22a_1
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3059_ _5071_/Q _5108_/Q VGND VGND VPWR VPWR _3059_/Y sky130_fd_sc_hd__nor2_1
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2430_ _2430_/A VGND VGND VPWR VPWR _2440_/B sky130_fd_sc_hd__inv_2
X_5080_ _3421_/X _5080_/D VGND VGND VPWR VPWR _5080_/Q sky130_fd_sc_hd__dfxtp_1
X_4100_ _4866_/Q _4099_/B _4099_/Y VGND VGND VPWR VPWR _4101_/A sky130_fd_sc_hd__a21oi_2
X_4031_ _4162_/A _4031_/B VGND VGND VPWR VPWR _4032_/B sky130_fd_sc_hd__or2_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4933_ _5047_/CLK _4933_/D VGND VGND VPWR VPWR _4933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ _5018_/CLK _4864_/D VGND VGND VPWR VPWR _4864_/Q sky130_fd_sc_hd__dfxtp_1
X_4795_ _2536_/X _4795_/D VGND VGND VPWR VPWR _4795_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3815_ _3815_/A VGND VGND VPWR VPWR _3817_/A sky130_fd_sc_hd__inv_2
X_3746_ _4935_/Q _3746_/B VGND VGND VPWR VPWR _3746_/Y sky130_fd_sc_hd__nor2_1
X_3677_ _3679_/A _3677_/B VGND VGND VPWR VPWR _5002_/D sky130_fd_sc_hd__nor2_1
X_2628_ _2628_/A VGND VGND VPWR VPWR _2774_/A sky130_fd_sc_hd__inv_2
X_2559_ _4737_/A _4733_/A _3318_/C _2554_/X VGND VGND VPWR VPWR _4790_/D sky130_fd_sc_hd__o211a_1
X_4229_ _4269_/A VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput11 dec_rate[4] VGND VGND VPWR VPWR _3532_/A sky130_fd_sc_hd__clkbuf_4
X_3600_ _3612_/A VGND VGND VPWR VPWR _3611_/A sky130_fd_sc_hd__clkbuf_2
X_4580_ _4580_/A VGND VGND VPWR VPWR _4587_/A sky130_fd_sc_hd__inv_2
X_3531_ _3531_/A _3531_/B _3531_/C VGND VGND VPWR VPWR _3531_/X sky130_fd_sc_hd__or3_1
X_3462_ _3978_/A VGND VGND VPWR VPWR _3462_/X sky130_fd_sc_hd__buf_2
X_3393_ _5090_/Q _3392_/Y _3375_/X _3393_/C1 VGND VGND VPWR VPWR _5090_/D sky130_fd_sc_hd__o211a_1
X_2413_ _2413_/A VGND VGND VPWR VPWR _2413_/Y sky130_fd_sc_hd__inv_2
X_5132_ _3176_/X _5132_/D VGND VGND VPWR VPWR _5132_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5063_ _5063_/CLK _5063_/D VGND VGND VPWR VPWR _5063_/Q sky130_fd_sc_hd__dfxtp_1
X_4014_ _4014_/A VGND VGND VPWR VPWR _4014_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4916_ _5028_/CLK _4916_/D VGND VGND VPWR VPWR _4916_/Q sky130_fd_sc_hd__dfxtp_1
X_4847_ _5028_/CLK _4847_/D VGND VGND VPWR VPWR _4847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4778_ _5047_/CLK _4778_/D VGND VGND VPWR VPWR _4778_/Q sky130_fd_sc_hd__dfxtp_1
X_3729_ _4868_/Q VGND VGND VPWR VPWR _4090_/A sky130_fd_sc_hd__inv_2
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2962_ _5095_/Q _5132_/Q VGND VGND VPWR VPWR _2962_/Y sky130_fd_sc_hd__nor2_1
X_4701_ _4631_/B _3029_/Y _4364_/X _5114_/Q VGND VGND VPWR VPWR _4702_/A sky130_fd_sc_hd__o22a_1
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4632_ _4632_/A _4632_/B VGND VGND VPWR VPWR _4838_/D sky130_fd_sc_hd__nor2_1
X_2893_ _5053_/Q VGND VGND VPWR VPWR _3478_/A sky130_fd_sc_hd__inv_2
XFILLER_8_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4563_ _4561_/Y _4550_/A _4562_/X _4557_/X VGND VGND VPWR VPWR _4875_/D sky130_fd_sc_hd__o211a_1
X_4494_ _4494_/A VGND VGND VPWR VPWR _4494_/Y sky130_fd_sc_hd__inv_2
X_3514_ _2864_/Y _3513_/A input3/X _3513_/Y VGND VGND VPWR VPWR _3514_/X sky130_fd_sc_hd__o22a_1
X_3445_ _3455_/A VGND VGND VPWR VPWR _3445_/X sky130_fd_sc_hd__buf_1
X_3376_ _5096_/Q _3374_/Y _3375_/X _3376_/C1 VGND VGND VPWR VPWR _5096_/D sky130_fd_sc_hd__o211a_1
X_5115_ _3261_/X _5115_/D VGND VGND VPWR VPWR _5115_/Q sky130_fd_sc_hd__dfxtp_1
X_5046_ _5047_/CLK _5046_/D VGND VGND VPWR VPWR _5046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3001_/A _3229_/Y _2996_/A _3229_/A _3193_/X VGND VGND VPWR VPWR _5122_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3161_ _2934_/Y _3160_/Y _2934_/A _3160_/A _3660_/A VGND VGND VPWR VPWR _5136_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3092_ _5064_/Q VGND VGND VPWR VPWR _3324_/A sky130_fd_sc_hd__clkinv_1
XFILLER_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3994_ _3994_/A _3994_/B VGND VGND VPWR VPWR _3995_/A sky130_fd_sc_hd__nand2_1
X_2945_ _2945_/A VGND VGND VPWR VPWR _2945_/X sky130_fd_sc_hd__clkbuf_2
X_2876_ input6/X _3498_/B _3494_/B VGND VGND VPWR VPWR _2876_/X sky130_fd_sc_hd__a21bo_1
X_4615_ _4621_/A VGND VGND VPWR VPWR _4620_/A sky130_fd_sc_hd__buf_2
X_4546_ _4546_/A VGND VGND VPWR VPWR _4546_/Y sky130_fd_sc_hd__inv_2
X_4477_ _4606_/B _4860_/Q _4481_/B VGND VGND VPWR VPWR _4478_/A sky130_fd_sc_hd__o21ai_1
X_3428_ _5078_/Q _3427_/Y _3406_/X _3428_/C1 VGND VGND VPWR VPWR _5078_/D sky130_fd_sc_hd__o211a_1
X_3359_ _3936_/A VGND VGND VPWR VPWR _3359_/X sky130_fd_sc_hd__buf_2
XFILLER_57_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5029_ _5047_/CLK _5029_/D VGND VGND VPWR VPWR _5029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2730_ _2730_/A _2730_/B _2730_/C _2730_/D VGND VGND VPWR VPWR _2735_/B sky130_fd_sc_hd__or4_4
X_2661_ _4955_/Q VGND VGND VPWR VPWR _2768_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4400_ _4400_/A VGND VGND VPWR VPWR _4400_/Y sky130_fd_sc_hd__inv_2
X_2592_ input6/X input7/X _3506_/Y input5/X VGND VGND VPWR VPWR _2593_/C sky130_fd_sc_hd__or4_4
X_4331_ _4331_/A VGND VGND VPWR VPWR _4335_/A sky130_fd_sc_hd__inv_2
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4262_ _4091_/Y _4261_/Y _4097_/A VGND VGND VPWR VPWR _4262_/Y sky130_fd_sc_hd__o21ai_1
X_3213_ _3212_/Y _2983_/A _3186_/X _3207_/X VGND VGND VPWR VPWR _5125_/D sky130_fd_sc_hd__o211a_1
X_4193_ _4481_/A _4193_/B _4193_/C VGND VGND VPWR VPWR _4924_/D sky130_fd_sc_hd__and3_1
X_3144_ _3354_/A _2945_/X _2940_/Y _3355_/A _3143_/Y VGND VGND VPWR VPWR _3144_/X
+ sky130_fd_sc_hd__o32a_1
X_3075_ _5071_/Q VGND VGND VPWR VPWR _3329_/A sky130_fd_sc_hd__clkinv_1
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3977_ _3974_/A _3973_/Y _3974_/Y _3973_/A _3976_/X VGND VGND VPWR VPWR _4948_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2928_ _3225_/A VGND VGND VPWR VPWR _3172_/A sky130_fd_sc_hd__buf_1
X_2859_ _2859_/A VGND VGND VPWR VPWR _2922_/C sky130_fd_sc_hd__inv_2
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4529_ _4623_/B _4846_/Q _4528_/X VGND VGND VPWR VPWR _4530_/A sky130_fd_sc_hd__o21ai_1
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 dec_rate[2] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_4
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3900_ _3591_/B _5041_/Q _3899_/Y VGND VGND VPWR VPWR _3901_/A sky130_fd_sc_hd__o21ai_1
X_4880_ _5028_/CLK _4880_/D VGND VGND VPWR VPWR _4880_/Q sky130_fd_sc_hd__dfxtp_1
X_3831_ _3831_/A _3994_/B VGND VGND VPWR VPWR _3845_/C sky130_fd_sc_hd__nand2_1
X_3762_ _4931_/Q _3762_/B VGND VGND VPWR VPWR _3762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2713_ _2778_/A VGND VGND VPWR VPWR _2713_/X sky130_fd_sc_hd__buf_1
X_3693_ _3726_/A VGND VGND VPWR VPWR _3703_/A sky130_fd_sc_hd__clkbuf_2
X_2644_ _4952_/Q VGND VGND VPWR VPWR _2736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2575_ _2636_/B _2691_/B VGND VGND VPWR VPWR _2575_/X sky130_fd_sc_hd__or2_1
X_4314_ _4617_/B _4851_/Q _4312_/X _4313_/Y VGND VGND VPWR VPWR _4315_/A sky130_fd_sc_hd__o22a_1
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4245_ _4240_/A _4240_/B _4220_/X _4240_/Y VGND VGND VPWR VPWR _4910_/D sky130_fd_sc_hd__o211a_1
X_4176_ _4176_/A VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__clkbuf_2
X_3127_ _3127_/A VGND VGND VPWR VPWR _3129_/B sky130_fd_sc_hd__inv_2
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3058_ _3058_/A _3058_/B VGND VGND VPWR VPWR _3058_/X sky130_fd_sc_hd__or2_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4030_ _4030_/A VGND VGND VPWR VPWR _4031_/B sky130_fd_sc_hd__inv_2
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4932_ _5047_/CLK _4932_/D VGND VGND VPWR VPWR _4932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4863_ _5018_/CLK _4863_/D VGND VGND VPWR VPWR _4863_/Q sky130_fd_sc_hd__dfxtp_1
X_4794_ _2543_/X _4794_/D VGND VGND VPWR VPWR _4794_/Q sky130_fd_sc_hd__dfxtp_1
X_3814_ _3639_/B _5020_/Q _4909_/Q _3813_/Y VGND VGND VPWR VPWR _3815_/A sky130_fd_sc_hd__o22a_1
X_3745_ _5046_/Q VGND VGND VPWR VPWR _3746_/B sky130_fd_sc_hd__inv_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3676_ _4891_/Q VGND VGND VPWR VPWR _3677_/B sky130_fd_sc_hd__inv_2
X_2627_ _2632_/D _2632_/B _2627_/C _4955_/Q VGND VGND VPWR VPWR _2628_/A sky130_fd_sc_hd__or4b_4
X_2558_ _2560_/A VGND VGND VPWR VPWR _2558_/X sky130_fd_sc_hd__buf_1
X_2489_ _2497_/A VGND VGND VPWR VPWR _2489_/X sky130_fd_sc_hd__buf_1
X_4228_ _4228_/A VGND VGND VPWR VPWR _4228_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4159_ _4019_/Y _4158_/Y _4019_/A _4158_/A _4151_/X VGND VGND VPWR VPWR _4933_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 dec_rate[5] VGND VGND VPWR VPWR _3516_/A sky130_fd_sc_hd__buf_2
X_3530_ _2895_/Y _3529_/X _2895_/Y _3529_/X VGND VGND VPWR VPWR _3531_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3461_ _3461_/A VGND VGND VPWR VPWR _3466_/B sky130_fd_sc_hd__inv_2
X_3392_ _3392_/A VGND VGND VPWR VPWR _3392_/Y sky130_fd_sc_hd__clkinvlp_2
X_2412_ _4606_/B _2937_/X _2411_/X VGND VGND VPWR VPWR _2413_/A sky130_fd_sc_hd__o21ai_1
XFILLER_69_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5131_ _3184_/X _5131_/D VGND VGND VPWR VPWR _5131_/Q sky130_fd_sc_hd__dfxtp_1
X_5062_ _5063_/CLK _5062_/D VGND VGND VPWR VPWR _5062_/Q sky130_fd_sc_hd__dfxtp_1
X_4013_ _4898_/Q _4012_/B _4012_/Y VGND VGND VPWR VPWR _4014_/A sky130_fd_sc_hd__a21oi_2
XFILLER_52_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4915_ _5028_/CLK _4915_/D VGND VGND VPWR VPWR _4915_/Q sky130_fd_sc_hd__dfxtp_1
X_4846_ _5028_/CLK _4846_/D VGND VGND VPWR VPWR _4846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4777_ _5047_/CLK _4777_/D VGND VGND VPWR VPWR _4777_/Q sky130_fd_sc_hd__dfxtp_1
X_3728_ _3736_/A _3728_/B VGND VGND VPWR VPWR _4980_/D sky130_fd_sc_hd__nor2_1
X_3659_ _3668_/A _3659_/B VGND VGND VPWR VPWR _5011_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2961_ _5094_/Q _5131_/Q _3352_/A _2960_/X VGND VGND VPWR VPWR _3180_/A sky130_fd_sc_hd__o22a_1
X_4700_ _4700_/A _4700_/B VGND VGND VPWR VPWR _4706_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4631_ _4632_/A _4631_/B VGND VGND VPWR VPWR _4839_/D sky130_fd_sc_hd__nor2_1
X_2892_ _3517_/A _2848_/B _2882_/Y VGND VGND VPWR VPWR _2894_/A sky130_fd_sc_hd__a21oi_4
X_4562_ _4562_/A VGND VGND VPWR VPWR _4562_/X sky130_fd_sc_hd__clkbuf_2
X_4493_ _4611_/B _4856_/Q _4492_/Y VGND VGND VPWR VPWR _4494_/A sky130_fd_sc_hd__o21ai_1
X_3513_ _3513_/A VGND VGND VPWR VPWR _3513_/Y sky130_fd_sc_hd__inv_2
X_3444_ _3444_/A VGND VGND VPWR VPWR _3455_/A sky130_fd_sc_hd__buf_1
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3375_ _3375_/A VGND VGND VPWR VPWR _3375_/X sky130_fd_sc_hd__buf_2
X_5114_ _3263_/X _5114_/D VGND VGND VPWR VPWR _5114_/Q sky130_fd_sc_hd__dfxtp_1
X_5045_ _5047_/CLK _5045_/D VGND VGND VPWR VPWR _5045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4829_ _5139_/Q _4829_/D VGND VGND VPWR VPWR _4829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3160_ _3160_/A VGND VGND VPWR VPWR _3160_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3091_ _5102_/Q VGND VGND VPWR VPWR _3091_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3993_ _3989_/A _3989_/B _3978_/X _3989_/Y VGND VGND VPWR VPWR _4943_/D sky130_fd_sc_hd__o211a_1
XFILLER_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2944_ _5133_/Q VGND VGND VPWR VPWR _2945_/A sky130_fd_sc_hd__inv_2
X_2875_ _5061_/Q VGND VGND VPWR VPWR _3487_/A sky130_fd_sc_hd__inv_2
X_4614_ _4614_/A _4614_/B VGND VGND VPWR VPWR _4853_/D sky130_fd_sc_hd__nor2_1
X_4545_ _4445_/A _4544_/Y _4441_/A _4544_/A _4539_/X VGND VGND VPWR VPWR _4880_/D
+ sky130_fd_sc_hd__o221a_1
X_4476_ _4480_/A _4480_/B VGND VGND VPWR VPWR _4481_/B sky130_fd_sc_hd__or2_1
X_3427_ _3427_/A VGND VGND VPWR VPWR _3427_/Y sky130_fd_sc_hd__inv_2
X_3358_ _3358_/A VGND VGND VPWR VPWR _3358_/Y sky130_fd_sc_hd__inv_2
X_3289_ _3289_/A VGND VGND VPWR VPWR _3289_/X sky130_fd_sc_hd__buf_1
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5028_ _5028_/CLK _5028_/D VGND VGND VPWR VPWR _5028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2660_ _2811_/A _2606_/B _2659_/X VGND VGND VPWR VPWR _2665_/C sky130_fd_sc_hd__o21a_1
XFILLER_8_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2591_ _3503_/X input3/X _2858_/A _2866_/A VGND VGND VPWR VPWR _2646_/A sky130_fd_sc_hd__or4b_4
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4330_ _4327_/X _4328_/Y _4622_/B _4847_/Q VGND VGND VPWR VPWR _4331_/A sky130_fd_sc_hd__o22a_1
X_4261_ _4261_/A VGND VGND VPWR VPWR _4261_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3212_ _3212_/A VGND VGND VPWR VPWR _3212_/Y sky130_fd_sc_hd__inv_2
X_4192_ _4192_/A _4192_/B VGND VGND VPWR VPWR _4193_/C sky130_fd_sc_hd__nand2_1
X_3143_ _5134_/Q VGND VGND VPWR VPWR _3143_/Y sky130_fd_sc_hd__inv_2
X_3074_ _3074_/A VGND VGND VPWR VPWR _3074_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3976_ _4269_/A VGND VGND VPWR VPWR _3976_/X sky130_fd_sc_hd__buf_2
X_2927_ _2927_/A VGND VGND VPWR VPWR _3225_/A sky130_fd_sc_hd__buf_1
XFILLER_50_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2858_ _2858_/A _3507_/B VGND VGND VPWR VPWR _2859_/A sky130_fd_sc_hd__or2_2
X_2789_ _4962_/Q _2787_/X _2788_/X VGND VGND VPWR VPWR _2800_/A sky130_fd_sc_hd__o21a_1
XFILLER_2_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4528_ _4532_/A _4528_/B VGND VGND VPWR VPWR _4528_/X sky130_fd_sc_hd__or2_1
X_4459_ _4614_/B _4853_/Q _4616_/B _4852_/Q VGND VGND VPWR VPWR _4459_/X sky130_fd_sc_hd__a211o_1
XFILLER_58_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2926__1 _5139_/CLK VGND VGND VPWR VPWR _3458_/A sky130_fd_sc_hd__inv_2
XFILLER_49_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3830_ _3825_/A _5015_/Q _3825_/Y VGND VGND VPWR VPWR _3994_/B sky130_fd_sc_hd__a21oi_4
X_3761_ _5042_/Q VGND VGND VPWR VPWR _3762_/B sky130_fd_sc_hd__inv_2
X_2712_ _2777_/A VGND VGND VPWR VPWR _2712_/X sky130_fd_sc_hd__buf_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3692_ _3692_/A _3692_/B VGND VGND VPWR VPWR _4996_/D sky130_fd_sc_hd__nor2_1
X_2643_ _2643_/A _2691_/B VGND VGND VPWR VPWR _2643_/X sky130_fd_sc_hd__or2_1
X_2574_ _2831_/B VGND VGND VPWR VPWR _2691_/B sky130_fd_sc_hd__buf_1
X_4313_ _4851_/Q VGND VGND VPWR VPWR _4313_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4244_ _4243_/A _4242_/Y _4243_/Y _4242_/A _4229_/X VGND VGND VPWR VPWR _4911_/D
+ sky130_fd_sc_hd__o221a_1
X_4175_ _4175_/A VGND VGND VPWR VPWR _4175_/Y sky130_fd_sc_hd__inv_2
X_3126_ _5087_/Q _5124_/Q _2986_/Y VGND VGND VPWR VPWR _3127_/A sky130_fd_sc_hd__a21oi_2
X_3057_ _3057_/A _3281_/B VGND VGND VPWR VPWR _3058_/B sky130_fd_sc_hd__or2_1
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3959_ _3628_/B _5025_/Q _3958_/Y VGND VGND VPWR VPWR _3960_/A sky130_fd_sc_hd__o21ai_1
XFILLER_2_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4931_ _5047_/CLK _4931_/D VGND VGND VPWR VPWR _4931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4862_ _5047_/CLK _4862_/D VGND VGND VPWR VPWR _4862_/Q sky130_fd_sc_hd__dfxtp_1
X_3813_ _5020_/Q VGND VGND VPWR VPWR _3813_/Y sky130_fd_sc_hd__inv_2
X_4793_ _2546_/X _4793_/D VGND VGND VPWR VPWR _4793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3744_ _3744_/A VGND VGND VPWR VPWR _3744_/Y sky130_fd_sc_hd__inv_2
X_3675_ _3679_/A _3675_/B VGND VGND VPWR VPWR _5003_/D sky130_fd_sc_hd__nor2_1
X_2626_ _4943_/Q _4944_/Q _2626_/C VGND VGND VPWR VPWR _2632_/D sky130_fd_sc_hd__or3_1
X_2557_ _4731_/Y _2556_/Y _4731_/A _2556_/A _2495_/X VGND VGND VPWR VPWR _4791_/D
+ sky130_fd_sc_hd__o221a_1
X_2488_ _4687_/A _2487_/B _2486_/X _2487_/Y VGND VGND VPWR VPWR _4807_/D sky130_fd_sc_hd__o211a_1
X_4227_ _3710_/B _4988_/Q _4226_/Y VGND VGND VPWR VPWR _4228_/A sky130_fd_sc_hd__o21ai_1
X_4158_ _4158_/A VGND VGND VPWR VPWR _4158_/Y sky130_fd_sc_hd__inv_2
X_3109_ _3333_/A _3041_/X _3332_/A _3045_/X VGND VGND VPWR VPWR _3109_/X sky130_fd_sc_hd__a211o_1
X_4089_ _3728_/B _4980_/Q _3728_/B _4980_/Q VGND VGND VPWR VPWR _4252_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput13 dec_rate[6] VGND VGND VPWR VPWR _2891_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3460_ _4648_/A VGND VGND VPWR VPWR _3460_/X sky130_fd_sc_hd__buf_1
X_3391_ _3396_/A VGND VGND VPWR VPWR _3391_/X sky130_fd_sc_hd__buf_1
X_2411_ _2416_/A _4654_/Y VGND VGND VPWR VPWR _2411_/X sky130_fd_sc_hd__or2_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5130_ _3188_/X _5130_/D VGND VGND VPWR VPWR _5130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5061_ _5063_/CLK _5061_/D VGND VGND VPWR VPWR _5061_/Q sky130_fd_sc_hd__dfxtp_1
X_4012_ _4898_/Q _4012_/B VGND VGND VPWR VPWR _4012_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4914_ _5028_/CLK _4914_/D VGND VGND VPWR VPWR _4914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4845_ _5028_/CLK _4845_/D VGND VGND VPWR VPWR _4845_/Q sky130_fd_sc_hd__dfxtp_1
X_4776_ _5047_/CLK _4776_/D VGND VGND VPWR VPWR _4776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3727_ _4869_/Q VGND VGND VPWR VPWR _3728_/B sky130_fd_sc_hd__inv_2
X_3658_ _4900_/Q VGND VGND VPWR VPWR _3659_/B sky130_fd_sc_hd__inv_2
X_3589_ _3612_/A VGND VGND VPWR VPWR _3599_/A sky130_fd_sc_hd__clkbuf_2
X_2609_ _4958_/Q _4960_/Q _4959_/Q _4961_/Q VGND VGND VPWR VPWR _2621_/C sky130_fd_sc_hd__or4_4
XFILLER_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2960_ _2960_/A VGND VGND VPWR VPWR _2960_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2891_ _2891_/A VGND VGND VPWR VPWR _3517_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4630_ _4632_/A _4630_/B VGND VGND VPWR VPWR _4840_/D sky130_fd_sc_hd__nor2_1
X_4561_ _4561_/A VGND VGND VPWR VPWR _4561_/Y sky130_fd_sc_hd__inv_2
X_4492_ _4492_/A _4492_/B VGND VGND VPWR VPWR _4492_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3512_ _3512_/A _3512_/B VGND VGND VPWR VPWR _3513_/A sky130_fd_sc_hd__nand2_1
X_3443_ _3331_/A _3443_/A2 _3431_/X _3440_/Y VGND VGND VPWR VPWR _5073_/D sky130_fd_sc_hd__a211oi_1
X_5113_ _3269_/X _5113_/D VGND VGND VPWR VPWR _5113_/Q sky130_fd_sc_hd__dfxtp_1
X_3374_ _3374_/A VGND VGND VPWR VPWR _3374_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5044_ _5047_/CLK _5044_/D VGND VGND VPWR VPWR _5044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4828_ _5139_/Q _4828_/D VGND VGND VPWR VPWR _4828_/Q sky130_fd_sc_hd__dfxtp_1
X_4759_ _2701_/X _2691_/X _4770_/S VGND VGND VPWR VPWR _4776_/D sky130_fd_sc_hd__mux2_2
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3090_ _3324_/C VGND VGND VPWR VPWR _3090_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3992_ _3845_/A _3991_/Y _3822_/A _3991_/A _3976_/X VGND VGND VPWR VPWR _4944_/D
+ sky130_fd_sc_hd__o221a_1
X_2943_ _5096_/Q VGND VGND VPWR VPWR _3354_/A sky130_fd_sc_hd__clkinvlp_4
X_2874_ _3483_/A _2870_/Y _5060_/Q _2863_/Y _2873_/Y VGND VGND VPWR VPWR _2874_/Y
+ sky130_fd_sc_hd__o221ai_2
X_4613_ _4614_/A _4613_/B VGND VGND VPWR VPWR _4854_/D sky130_fd_sc_hd__nor2_1
X_4544_ _4544_/A VGND VGND VPWR VPWR _4544_/Y sky130_fd_sc_hd__inv_2
X_4475_ _4277_/Y _4474_/A _4277_/A _4474_/Y _4269_/X VGND VGND VPWR VPWR _4899_/D
+ sky130_fd_sc_hd__o221a_1
X_3426_ _3426_/A VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__buf_1
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3357_ _3357_/A _3357_/B VGND VGND VPWR VPWR _3358_/A sky130_fd_sc_hd__or2_4
X_3288_ _3286_/Y _3056_/A _3287_/X _3281_/X VGND VGND VPWR VPWR _5109_/D sky130_fd_sc_hd__o211a_1
X_5027_ _5028_/CLK _5027_/D VGND VGND VPWR VPWR _5027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ _2590_/A _2590_/B _2590_/C _2590_/D VGND VGND VPWR VPWR _2590_/X sky130_fd_sc_hd__or4_4
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4260_ _4260_/A _4260_/B VGND VGND VPWR VPWR _4261_/A sky130_fd_sc_hd__nand2_1
X_4191_ _4040_/A _4189_/Y _4038_/A _4189_/A _4190_/X VGND VGND VPWR VPWR _4925_/D
+ sky130_fd_sc_hd__o221a_1
X_3211_ _3222_/A VGND VGND VPWR VPWR _3211_/X sky130_fd_sc_hd__buf_1
XFILLER_79_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3142_ _5097_/Q VGND VGND VPWR VPWR _3355_/A sky130_fd_sc_hd__clkinv_1
X_3073_ _5069_/Q _5106_/Q _3069_/Y _3072_/Y VGND VGND VPWR VPWR _3074_/A sky130_fd_sc_hd__o22a_1
XFILLER_27_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3975_ _4500_/A VGND VGND VPWR VPWR _4269_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2857_ _2857_/A VGND VGND VPWR VPWR _3507_/B sky130_fd_sc_hd__buf_1
X_2788_ _2788_/A VGND VGND VPWR VPWR _2788_/X sky130_fd_sc_hd__buf_1
X_4527_ _4522_/A _4522_/B _4526_/X _4522_/Y VGND VGND VPWR VPWR _4885_/D sky130_fd_sc_hd__o211a_1
X_4458_ _4458_/A VGND VGND VPWR VPWR _4616_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_77_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3409_ _3343_/A _3409_/A2 _3401_/X _3404_/Y VGND VGND VPWR VPWR _5085_/D sky130_fd_sc_hd__a211oi_1
X_4389_ _4795_/Q _4389_/B VGND VGND VPWR VPWR _4389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2926__2 _5139_/CLK VGND VGND VPWR VPWR _3246_/A sky130_fd_sc_hd__inv_2
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3760_ _3591_/B _5041_/Q _3591_/B _5041_/Q VGND VGND VPWR VPWR _3895_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2711_ _4944_/Q _2709_/X _2710_/X VGND VGND VPWR VPWR _2715_/C sky130_fd_sc_hd__o21a_1
X_3691_ _3691_/A VGND VGND VPWR VPWR _3692_/B sky130_fd_sc_hd__buf_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2642_ _2658_/A _2606_/Y _2662_/A _2613_/Y _2641_/X VGND VGND VPWR VPWR _2642_/Y
+ sky130_fd_sc_hd__o221ai_1
X_2573_ _2632_/B _2573_/B _2603_/D _2627_/C VGND VGND VPWR VPWR _2831_/B sky130_fd_sc_hd__nor4_2
X_4312_ _4813_/Q VGND VGND VPWR VPWR _4312_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4243_ _4243_/A VGND VGND VPWR VPWR _4243_/Y sky130_fd_sc_hd__inv_2
X_4174_ _4025_/B _4173_/Y _4024_/A _4173_/A _4151_/X VGND VGND VPWR VPWR _4929_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3125_ _3125_/A _3125_/B VGND VGND VPWR VPWR _3129_/A sky130_fd_sc_hd__or2_1
XFILLER_67_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3056_ _3056_/A VGND VGND VPWR VPWR _3281_/B sky130_fd_sc_hd__inv_2
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3958_ _3958_/A _3958_/B VGND VGND VPWR VPWR _3958_/Y sky130_fd_sc_hd__nand2_1
X_3889_ _3893_/A _3893_/B VGND VGND VPWR VPWR _3894_/B sky130_fd_sc_hd__or2_1
X_2909_ _3525_/A _2908_/X _3525_/A _2908_/X VGND VGND VPWR VPWR _2914_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ _5047_/CLK _4930_/D VGND VGND VPWR VPWR _4930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4861_ _5047_/CLK _4861_/D VGND VGND VPWR VPWR _4861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3812_ _3974_/A _3969_/A VGND VGND VPWR VPWR _3818_/A sky130_fd_sc_hd__or2_1
X_4792_ _2551_/X _4792_/D VGND VGND VPWR VPWR _4792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3743_ _4936_/Q _5047_/Q _4936_/Q _5047_/Q VGND VGND VPWR VPWR _3744_/A sky130_fd_sc_hd__a2bb2o_1
X_3674_ _4892_/Q VGND VGND VPWR VPWR _3675_/B sky130_fd_sc_hd__inv_2
X_2625_ _4942_/Q _4939_/Q _4940_/Q _4941_/Q VGND VGND VPWR VPWR _2626_/C sky130_fd_sc_hd__or4_4
X_2556_ _2556_/A VGND VGND VPWR VPWR _2556_/Y sky130_fd_sc_hd__inv_2
X_2487_ _4687_/A _2487_/B VGND VGND VPWR VPWR _2487_/Y sky130_fd_sc_hd__nand2_1
X_4226_ _4226_/A _4226_/B VGND VGND VPWR VPWR _4226_/Y sky130_fd_sc_hd__nand2_1
X_4157_ _3668_/B _5006_/Q _4161_/B VGND VGND VPWR VPWR _4158_/A sky130_fd_sc_hd__o21ai_1
X_3108_ _5073_/Q _3050_/X _3107_/X VGND VGND VPWR VPWR _3108_/Y sky130_fd_sc_hd__o21ai_1
X_4088_ _4088_/A VGND VGND VPWR VPWR _4111_/A sky130_fd_sc_hd__inv_2
X_3039_ _5075_/Q VGND VGND VPWR VPWR _3333_/A sky130_fd_sc_hd__inv_1
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput14 dec_rate[7] VGND VGND VPWR VPWR _2881_/A sky130_fd_sc_hd__buf_1
XFILLER_10_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2410_ _2428_/A VGND VGND VPWR VPWR _2410_/X sky130_fd_sc_hd__buf_1
X_3390_ _3349_/A _3390_/A2 _3371_/X _3387_/Y VGND VGND VPWR VPWR _5091_/D sky130_fd_sc_hd__a211oi_1
X_5060_ _5063_/CLK _5060_/D VGND VGND VPWR VPWR _5060_/Q sky130_fd_sc_hd__dfxtp_2
X_4011_ _5009_/Q VGND VGND VPWR VPWR _4012_/B sky130_fd_sc_hd__inv_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4913_ _5028_/CLK _4913_/D VGND VGND VPWR VPWR _4913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4844_ _5028_/CLK _4844_/D VGND VGND VPWR VPWR _4844_/Q sky130_fd_sc_hd__dfxtp_1
X_4775_ _5018_/CLK _4775_/D VGND VGND VPWR VPWR _4775_/Q sky130_fd_sc_hd__dfxtp_1
X_3726_ _3726_/A VGND VGND VPWR VPWR _3736_/A sky130_fd_sc_hd__clkbuf_2
X_3657_ _3669_/A VGND VGND VPWR VPWR _3668_/A sky130_fd_sc_hd__buf_2
X_3588_ _3588_/A _3588_/B VGND VGND VPWR VPWR _5042_/D sky130_fd_sc_hd__nor2_1
X_2608_ _4956_/Q _4955_/Q _4954_/Q _4957_/Q VGND VGND VPWR VPWR _2620_/D sky130_fd_sc_hd__or4_4
X_2539_ _4720_/A _2539_/B VGND VGND VPWR VPWR _2539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4209_ _4219_/A _4127_/B _4056_/Y VGND VGND VPWR VPWR _4210_/B sky130_fd_sc_hd__o21ai_1
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2890_ _5055_/Q VGND VGND VPWR VPWR _3480_/A sky130_fd_sc_hd__inv_2
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4560_ _4371_/A _4559_/Y _4367_/A _4559_/A _4539_/X VGND VGND VPWR VPWR _4876_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4491_ _4305_/A _4497_/B _4454_/Y VGND VGND VPWR VPWR _4492_/B sky130_fd_sc_hd__o21ai_1
X_3511_ _3518_/A VGND VGND VPWR VPWR _3512_/A sky130_fd_sc_hd__inv_2
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3442_ _3442_/A VGND VGND VPWR VPWR _3442_/X sky130_fd_sc_hd__buf_1
X_3373_ _3382_/A VGND VGND VPWR VPWR _3373_/X sky130_fd_sc_hd__buf_1
X_5112_ _3272_/X _5112_/D VGND VGND VPWR VPWR _5112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5043_ _5047_/CLK _5043_/D VGND VGND VPWR VPWR _5043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _5018_/CLK _4827_/D VGND VGND VPWR VPWR _4827_/Q sky130_fd_sc_hd__dfxtp_1
X_4758_ _2690_/X _2680_/X _4770_/S VGND VGND VPWR VPWR _4775_/D sky130_fd_sc_hd__mux2_1
X_4689_ _4343_/X _3011_/X _4688_/X VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__o21ai_1
X_3709_ _4877_/Q VGND VGND VPWR VPWR _3710_/B sky130_fd_sc_hd__inv_2
XFILLER_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3991_ _3991_/A VGND VGND VPWR VPWR _3991_/Y sky130_fd_sc_hd__inv_2
X_2942_ _2942_/A VGND VGND VPWR VPWR _2942_/Y sky130_fd_sc_hd__inv_2
X_2873_ _3481_/A _2872_/Y _3483_/A _2870_/Y VGND VGND VPWR VPWR _2873_/Y sky130_fd_sc_hd__a22oi_2
X_4612_ _4614_/A _4612_/B VGND VGND VPWR VPWR _4855_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4543_ _4628_/B _4842_/Q _4542_/X VGND VGND VPWR VPWR _4544_/A sky130_fd_sc_hd__o21ai_1
X_4474_ _4474_/A VGND VGND VPWR VPWR _4474_/Y sky130_fd_sc_hd__inv_2
X_3425_ _3337_/A _3425_/A2 _3401_/X _3422_/Y VGND VGND VPWR VPWR _5079_/D sky130_fd_sc_hd__a211oi_1
X_3356_ _3356_/A _3356_/B VGND VGND VPWR VPWR _3357_/B sky130_fd_sc_hd__or2_2
X_3287_ _3375_/A VGND VGND VPWR VPWR _3287_/X sky130_fd_sc_hd__buf_2
XFILLER_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5026_ _5028_/CLK _5026_/D VGND VGND VPWR VPWR _5026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3210_ _2984_/A _3209_/Y _2979_/A _3209_/A _3193_/X VGND VGND VPWR VPWR _5126_/D
+ sky130_fd_sc_hd__o221a_1
X_4190_ _4269_/A VGND VGND VPWR VPWR _4190_/X sky130_fd_sc_hd__buf_2
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3141_ _2965_/X _2985_/X _3212_/A _3140_/X VGND VGND VPWR VPWR _3173_/A sky130_fd_sc_hd__o31a_1
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3072_ _3326_/A _4722_/B VGND VGND VPWR VPWR _3072_/Y sky130_fd_sc_hd__nor2_4
XFILLER_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3974_ _3974_/A VGND VGND VPWR VPWR _3974_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2925_ _5138_/Q _2842_/Y _4771_/X _4647_/B _3612_/A VGND VGND VPWR VPWR _5138_/D
+ sky130_fd_sc_hd__a221o_1
X_2856_ input6/X input7/X input4/X input5/X VGND VGND VPWR VPWR _2858_/A sky130_fd_sc_hd__or4_4
X_2787_ _2787_/A VGND VGND VPWR VPWR _2787_/X sky130_fd_sc_hd__buf_1
X_4526_ _4562_/A VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__clkbuf_2
X_4457_ _4312_/X _4313_/Y _4456_/Y VGND VGND VPWR VPWR _4457_/Y sky130_fd_sc_hd__o21ai_1
X_3408_ _3413_/A VGND VGND VPWR VPWR _3408_/X sky130_fd_sc_hd__buf_1
X_4388_ _4833_/Q VGND VGND VPWR VPWR _4389_/B sky130_fd_sc_hd__inv_2
X_3339_ _3339_/A _3339_/B VGND VGND VPWR VPWR _3340_/B sky130_fd_sc_hd__or2_1
X_5009_ _5047_/CLK _5009_/D VGND VGND VPWR VPWR _5009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2926__3 _5139_/CLK VGND VGND VPWR VPWR _2927_/A sky130_fd_sc_hd__inv_2
XFILLER_64_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2710_ _2775_/A VGND VGND VPWR VPWR _2710_/X sky130_fd_sc_hd__buf_1
X_3690_ _4885_/Q VGND VGND VPWR VPWR _3691_/A sky130_fd_sc_hd__inv_2
X_2641_ _2646_/A _2617_/Y _2588_/A _2624_/Y _2640_/X VGND VGND VPWR VPWR _2641_/X
+ sky130_fd_sc_hd__o221a_1
X_2572_ _2616_/A _2631_/A VGND VGND VPWR VPWR _2627_/C sky130_fd_sc_hd__or2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4311_ _4813_/Q VGND VGND VPWR VPWR _4617_/B sky130_fd_sc_hd__inv_2
X_4242_ _4242_/A VGND VGND VPWR VPWR _4242_/Y sky130_fd_sc_hd__inv_2
X_4173_ _4173_/A VGND VGND VPWR VPWR _4173_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3124_ _3124_/A _3242_/B VGND VGND VPWR VPWR _3125_/B sky130_fd_sc_hd__or2_1
X_3055_ _3330_/A _3054_/Y _5072_/Q _5109_/Q VGND VGND VPWR VPWR _3056_/A sky130_fd_sc_hd__o22a_1
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3957_ _3809_/B _3963_/B _3848_/Y VGND VGND VPWR VPWR _3958_/B sky130_fd_sc_hd__o21ai_1
X_2908_ _3532_/A _2846_/B _2907_/Y VGND VGND VPWR VPWR _2908_/X sky130_fd_sc_hd__a21o_1
X_3888_ _3985_/A _3888_/B _3888_/C VGND VGND VPWR VPWR _4971_/D sky130_fd_sc_hd__and3_1
X_2839_ _4969_/Q _2783_/A _2798_/X VGND VGND VPWR VPWR _2840_/D sky130_fd_sc_hd__o21a_1
X_4509_ _4509_/A VGND VGND VPWR VPWR _4509_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4860_ _5047_/CLK _4860_/D VGND VGND VPWR VPWR _4860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3811_ _3637_/B _5021_/Q _3637_/B _5021_/Q VGND VGND VPWR VPWR _3969_/A sky130_fd_sc_hd__a2bb2o_1
X_4791_ _2553_/X _4791_/D VGND VGND VPWR VPWR _4791_/Q sky130_fd_sc_hd__dfxtp_2
X_3742_ _4601_/A _3742_/B VGND VGND VPWR VPWR _4974_/D sky130_fd_sc_hd__nor2_1
X_3673_ _3679_/A _3673_/B VGND VGND VPWR VPWR _5004_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2624_ _2680_/A _2624_/B VGND VGND VPWR VPWR _2624_/Y sky130_fd_sc_hd__nor2_1
X_2555_ _4644_/B _3086_/X _2554_/X VGND VGND VPWR VPWR _2556_/A sky130_fd_sc_hd__o21ai_1
X_2486_ _3165_/A VGND VGND VPWR VPWR _2486_/X sky130_fd_sc_hd__clkbuf_2
X_4225_ _4075_/B _4232_/B _4114_/Y VGND VGND VPWR VPWR _4226_/B sky130_fd_sc_hd__o21ai_1
X_4156_ _4160_/A _4160_/B VGND VGND VPWR VPWR _4161_/B sky130_fd_sc_hd__or2_1
X_3107_ _5073_/Q _3050_/X _5072_/Q _5109_/Q VGND VGND VPWR VPWR _3107_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4087_ _4870_/Q _4086_/B _4086_/Y VGND VGND VPWR VPWR _4088_/A sky130_fd_sc_hd__a21oi_2
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3038_ _3038_/A _3038_/B VGND VGND VPWR VPWR _3038_/X sky130_fd_sc_hd__or2_1
XFILLER_62_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4989_ _5028_/CLK _4989_/D VGND VGND VPWR VPWR _4989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 dec_rate[8] VGND VGND VPWR VPWR _2850_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4010_ _4010_/A VGND VGND VPWR VPWR _4010_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4912_ _5028_/CLK _4912_/D VGND VGND VPWR VPWR _4912_/Q sky130_fd_sc_hd__dfxtp_1
X_4843_ _5028_/CLK _4843_/D VGND VGND VPWR VPWR _4843_/Q sky130_fd_sc_hd__dfxtp_1
X_4774_ _5018_/CLK _4774_/D VGND VGND VPWR VPWR _4774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3725_ _3725_/A _3725_/B VGND VGND VPWR VPWR _4981_/D sky130_fd_sc_hd__nor2_1
X_3656_ _3656_/A _3656_/B VGND VGND VPWR VPWR _5012_/D sky130_fd_sc_hd__nor2_1
X_3587_ _4931_/Q VGND VGND VPWR VPWR _3588_/B sky130_fd_sc_hd__inv_2
X_2607_ _4954_/Q VGND VGND VPWR VPWR _2756_/A sky130_fd_sc_hd__clkbuf_2
X_2538_ _4728_/A _4728_/B _2547_/A _4724_/A VGND VGND VPWR VPWR _2539_/B sky130_fd_sc_hd__a31o_1
XFILLER_75_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2469_ _4620_/B _2991_/X _2468_/Y VGND VGND VPWR VPWR _2470_/A sky130_fd_sc_hd__o21ai_1
X_4208_ _4208_/A VGND VGND VPWR VPWR _4210_/A sky130_fd_sc_hd__inv_2
XFILLER_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4139_ _3673_/B _5004_/Q _4028_/Y _3671_/B _5005_/Q VGND VGND VPWR VPWR _4139_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3510_ _5060_/Q _3509_/X _5060_/Q _3509_/X VGND VGND VPWR VPWR _3544_/B sky130_fd_sc_hd__a2bb2o_1
X_4490_ _4490_/A VGND VGND VPWR VPWR _4497_/B sky130_fd_sc_hd__inv_2
X_3441_ _5074_/Q _3440_/Y _3435_/X _3441_/C1 VGND VGND VPWR VPWR _5074_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3372_ _3355_/A _3376_/C1 _3371_/X _3366_/Y VGND VGND VPWR VPWR _5097_/D sky130_fd_sc_hd__a211oi_1
XFILLER_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5111_ _3278_/X _5111_/D VGND VGND VPWR VPWR _5111_/Q sky130_fd_sc_hd__dfxtp_1
X_5042_ _5047_/CLK _5042_/D VGND VGND VPWR VPWR _5042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4826_ _5018_/CLK _4826_/D VGND VGND VPWR VPWR _4826_/Q sky130_fd_sc_hd__dfxtp_1
X_4757_ _2679_/X _2666_/X _4770_/S VGND VGND VPWR VPWR _4774_/D sky130_fd_sc_hd__mux2_1
X_4688_ _4343_/X _5118_/Q _4804_/Q _5117_/Q VGND VGND VPWR VPWR _4688_/X sky130_fd_sc_hd__a22o_1
X_3708_ _3714_/A _3708_/B VGND VGND VPWR VPWR _4989_/D sky130_fd_sc_hd__nor2_1
X_3639_ _3645_/A _3639_/B VGND VGND VPWR VPWR _5020_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3990_ _3645_/B _5017_/Q _3989_/Y VGND VGND VPWR VPWR _3991_/A sky130_fd_sc_hd__o21ai_1
X_2941_ _5097_/Q _5134_/Q _2940_/Y VGND VGND VPWR VPWR _2942_/A sky130_fd_sc_hd__a21oi_2
X_4611_ _4614_/A _4611_/B VGND VGND VPWR VPWR _4856_/D sky130_fd_sc_hd__nor2_1
X_2872_ _3501_/A _3502_/B _3503_/B VGND VGND VPWR VPWR _2872_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_30_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4542_ _4546_/A _4542_/B VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__or2_1
X_4473_ _4281_/Y _4480_/B _4480_/A _4472_/X VGND VGND VPWR VPWR _4474_/A sky130_fd_sc_hd__o31a_1
XFILLER_7_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3424_ _3426_/A VGND VGND VPWR VPWR _3424_/X sky130_fd_sc_hd__buf_1
X_3355_ _3355_/A _3355_/B VGND VGND VPWR VPWR _3356_/B sky130_fd_sc_hd__or2_1
X_3286_ _3286_/A VGND VGND VPWR VPWR _3286_/Y sky130_fd_sc_hd__inv_2
X_5025_ _5028_/CLK _5025_/D VGND VGND VPWR VPWR _5025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4809_ _2474_/X _4809_/D VGND VGND VPWR VPWR _4809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3140_ _2965_/B _3132_/Y _2965_/X _3136_/X _3139_/X VGND VGND VPWR VPWR _3140_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3071_ _5105_/Q VGND VGND VPWR VPWR _4722_/B sky130_fd_sc_hd__clkinv_4
XFILLER_35_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3973_ _3973_/A VGND VGND VPWR VPWR _3973_/Y sky130_fd_sc_hd__inv_2
X_2924_ _3370_/A VGND VGND VPWR VPWR _3612_/A sky130_fd_sc_hd__clkbuf_4
X_2855_ input6/X _3498_/B VGND VGND VPWR VPWR _3494_/B sky130_fd_sc_hd__or2_2
X_2786_ _2786_/A _2821_/B VGND VGND VPWR VPWR _2786_/X sky130_fd_sc_hd__or2_1
X_4525_ _4450_/B _4524_/Y _4448_/A _4524_/A _4501_/X VGND VGND VPWR VPWR _4886_/D
+ sky130_fd_sc_hd__o221a_1
X_4456_ _4617_/B _4851_/Q _4618_/B _4850_/Q VGND VGND VPWR VPWR _4456_/Y sky130_fd_sc_hd__o22ai_1
X_3407_ _5086_/Q _3404_/Y _3406_/X _3407_/C1 VGND VGND VPWR VPWR _5086_/D sky130_fd_sc_hd__o211a_1
X_4387_ _4387_/A _4387_/B VGND VGND VPWR VPWR _4387_/X sky130_fd_sc_hd__or2_1
XFILLER_49_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3338_ _3338_/A _3338_/B VGND VGND VPWR VPWR _3339_/B sky130_fd_sc_hd__or2_1
X_3269_ _3269_/A VGND VGND VPWR VPWR _3269_/X sky130_fd_sc_hd__buf_1
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5008_ _5047_/CLK _5008_/D VGND VGND VPWR VPWR _5008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2640_ _2585_/A _2630_/Y _2582_/A _2650_/A _2639_/Y VGND VGND VPWR VPWR _2640_/X
+ sky130_fd_sc_hd__o221a_1
X_2571_ _4946_/Q _4945_/Q _4948_/Q _4947_/Q VGND VGND VPWR VPWR _2631_/A sky130_fd_sc_hd__or4_4
X_4310_ _4510_/A _4505_/A VGND VGND VPWR VPWR _4320_/A sky130_fd_sc_hd__or2_1
X_4241_ _3719_/B _4984_/Q _4240_/Y VGND VGND VPWR VPWR _4242_/A sky130_fd_sc_hd__o21ai_1
X_4172_ _3677_/B _5002_/Q _4171_/X VGND VGND VPWR VPWR _4173_/A sky130_fd_sc_hd__o21ai_1
X_3123_ _3123_/A VGND VGND VPWR VPWR _3242_/B sky130_fd_sc_hd__inv_2
XFILLER_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3054_ _5109_/Q VGND VGND VPWR VPWR _3054_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3956_ _3956_/A VGND VGND VPWR VPWR _3963_/B sky130_fd_sc_hd__inv_2
X_2907_ _3515_/B VGND VGND VPWR VPWR _2907_/Y sky130_fd_sc_hd__inv_2
X_3887_ _3887_/A _3887_/B VGND VGND VPWR VPWR _3888_/C sky130_fd_sc_hd__nand2_1
X_2838_ _4972_/Q _2781_/A _2796_/X VGND VGND VPWR VPWR _2840_/C sky130_fd_sc_hd__o21a_1
X_2769_ _2567_/X _2722_/X _2723_/X VGND VGND VPWR VPWR _2785_/A sky130_fd_sc_hd__o21a_1
X_4508_ _4616_/B _4852_/Q _4507_/Y VGND VGND VPWR VPWR _4509_/A sky130_fd_sc_hd__o21ai_1
X_4439_ _4805_/Q VGND VGND VPWR VPWR _4626_/B sky130_fd_sc_hd__inv_2
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4790_ _2558_/X _4790_/D VGND VGND VPWR VPWR _4790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3810_ _3634_/B _5022_/Q _3634_/B _5022_/Q VGND VGND VPWR VPWR _3974_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3741_ _4863_/Q VGND VGND VPWR VPWR _3742_/B sky130_fd_sc_hd__inv_2
XFILLER_9_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ _4893_/Q VGND VGND VPWR VPWR _3673_/B sky130_fd_sc_hd__inv_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2623_ _2777_/A VGND VGND VPWR VPWR _2624_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2554_ _4737_/Y _4733_/Y VGND VGND VPWR VPWR _2554_/X sky130_fd_sc_hd__or2_1
X_2485_ _4625_/B _3008_/X _2484_/Y VGND VGND VPWR VPWR _2487_/B sky130_fd_sc_hd__o21ai_1
X_4224_ _4224_/A VGND VGND VPWR VPWR _4232_/B sky130_fd_sc_hd__inv_2
X_4155_ _4481_/A _4155_/B _4155_/C VGND VGND VPWR VPWR _4934_/D sky130_fd_sc_hd__and3_1
X_3106_ _5077_/Q _3030_/X _3105_/X VGND VGND VPWR VPWR _3106_/Y sky130_fd_sc_hd__o21ai_1
X_4086_ _4870_/Q _4086_/B VGND VGND VPWR VPWR _4086_/Y sky130_fd_sc_hd__nor2_1
X_3037_ _3037_/A _3264_/A VGND VGND VPWR VPWR _3038_/B sky130_fd_sc_hd__or2_1
XFILLER_36_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4988_ _5028_/CLK _4988_/D VGND VGND VPWR VPWR _4988_/Q sky130_fd_sc_hd__dfxtp_1
X_3939_ _3978_/A VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput16 dec_rate[9] VGND VGND VPWR VPWR _3501_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4911_ _5028_/CLK _4911_/D VGND VGND VPWR VPWR _4911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4842_ _5028_/CLK _4842_/D VGND VGND VPWR VPWR _4842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4773_ _5018_/CLK _4773_/D VGND VGND VPWR VPWR _4773_/Q sky130_fd_sc_hd__dfxtp_1
X_3724_ _4870_/Q VGND VGND VPWR VPWR _3725_/B sky130_fd_sc_hd__inv_2
X_3655_ _4901_/Q VGND VGND VPWR VPWR _3656_/B sky130_fd_sc_hd__inv_2
X_2606_ _2801_/A _2606_/B VGND VGND VPWR VPWR _2606_/Y sky130_fd_sc_hd__nor2_1
X_3586_ _3588_/A _3586_/B VGND VGND VPWR VPWR _5043_/D sky130_fd_sc_hd__nor2_1
X_2537_ _4740_/D VGND VGND VPWR VPWR _2547_/A sky130_fd_sc_hd__inv_2
X_2468_ _2468_/A _2468_/B VGND VGND VPWR VPWR _2468_/Y sky130_fd_sc_hd__nand2_1
X_4207_ _4206_/Y _4195_/A _4177_/X _4202_/X VGND VGND VPWR VPWR _4920_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2399_ _4611_/B _2960_/X _4666_/Y _4610_/B _3138_/Y VGND VGND VPWR VPWR _2399_/X
+ sky130_fd_sc_hd__o32a_1
X_4138_ _3679_/B _5001_/Q _4041_/A _4136_/Y _4137_/X VGND VGND VPWR VPWR _4138_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4069_ _4069_/A _4222_/A VGND VGND VPWR VPWR _4075_/A sky130_fd_sc_hd__or2_1
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3440_ _3440_/A VGND VGND VPWR VPWR _3440_/Y sky130_fd_sc_hd__inv_2
X_3371_ _4639_/A VGND VGND VPWR VPWR _3371_/X sky130_fd_sc_hd__buf_2
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5110_ _3280_/X _5110_/D VGND VGND VPWR VPWR _5110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5041_ _5047_/CLK _5041_/D VGND VGND VPWR VPWR _5041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4825_ _5139_/CLK _4825_/D VGND VGND VPWR VPWR _4825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4756_ _2665_/X _2643_/X _4770_/S VGND VGND VPWR VPWR _4773_/D sky130_fd_sc_hd__mux2_1
X_4687_ _4687_/A _4687_/B VGND VGND VPWR VPWR _4687_/Y sky130_fd_sc_hd__nand2_1
X_3707_ _4878_/Q VGND VGND VPWR VPWR _3708_/B sky130_fd_sc_hd__inv_2
X_3638_ _4909_/Q VGND VGND VPWR VPWR _3639_/B sky130_fd_sc_hd__inv_2
X_3569_ _5054_/Q _3568_/Y _3480_/B _3559_/X VGND VGND VPWR VPWR _5054_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2940_ _5097_/Q _5134_/Q VGND VGND VPWR VPWR _2940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2871_ _5056_/Q VGND VGND VPWR VPWR _3481_/A sky130_fd_sc_hd__clkbuf_2
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4610_ _4614_/A _4610_/B VGND VGND VPWR VPWR _4857_/D sky130_fd_sc_hd__nor2_1
X_4541_ _4536_/A _4536_/B _4526_/X _4536_/Y VGND VGND VPWR VPWR _4881_/D sky130_fd_sc_hd__o211a_1
X_4472_ _4606_/B _4860_/Q _4279_/Y _4605_/B _4861_/Q VGND VGND VPWR VPWR _4472_/X
+ sky130_fd_sc_hd__o32a_1
X_3423_ _5080_/Q _3422_/Y _3406_/X _3423_/C1 VGND VGND VPWR VPWR _5080_/D sky130_fd_sc_hd__o211a_1
X_3354_ _3354_/A _3354_/B VGND VGND VPWR VPWR _3355_/B sky130_fd_sc_hd__or2_1
X_3285_ _3289_/A VGND VGND VPWR VPWR _3285_/X sky130_fd_sc_hd__buf_1
X_5024_ _5028_/CLK _5024_/D VGND VGND VPWR VPWR _5024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4808_ _2480_/X _4808_/D VGND VGND VPWR VPWR _4808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4739_ _4731_/Y _4733_/Y _4737_/Y _4738_/X VGND VGND VPWR VPWR _4740_/D sky130_fd_sc_hd__o31a_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3070_ _5068_/Q VGND VGND VPWR VPWR _3326_/A sky130_fd_sc_hd__inv_2
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3972_ _3637_/B _5021_/Q _3971_/Y VGND VGND VPWR VPWR _3973_/A sky130_fd_sc_hd__o21ai_1
X_2923_ _5138_/Q _2923_/B VGND VGND VPWR VPWR _4647_/B sky130_fd_sc_hd__nand2_1
X_2854_ input5/X _3508_/B VGND VGND VPWR VPWR _3498_/B sky130_fd_sc_hd__or2_1
X_2785_ _2785_/A _2785_/B _2785_/C _2785_/D VGND VGND VPWR VPWR _2785_/X sky130_fd_sc_hd__or4_1
X_4524_ _4524_/A VGND VGND VPWR VPWR _4524_/Y sky130_fd_sc_hd__inv_2
X_4455_ _4455_/A VGND VGND VPWR VPWR _4614_/B sky130_fd_sc_hd__clkbuf_2
X_3406_ _3978_/A VGND VGND VPWR VPWR _3406_/X sky130_fd_sc_hd__clkbuf_2
X_4386_ _4386_/A _4577_/B VGND VGND VPWR VPWR _4387_/B sky130_fd_sc_hd__or2_1
X_3337_ _3337_/A _3337_/B VGND VGND VPWR VPWR _3338_/B sky130_fd_sc_hd__or2_1
XFILLER_58_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3268_ _3037_/A _3266_/Y _3032_/A _3266_/A _3267_/X VGND VGND VPWR VPWR _5114_/D
+ sky130_fd_sc_hd__o221a_1
X_5007_ _5047_/CLK _5007_/D VGND VGND VPWR VPWR _5007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3199_ _3199_/A _3199_/B VGND VGND VPWR VPWR _3199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2570_ _4951_/Q _4952_/Q _4954_/Q _4953_/Q VGND VGND VPWR VPWR _2616_/A sky130_fd_sc_hd__or4_4
X_4240_ _4240_/A _4240_/B VGND VGND VPWR VPWR _4240_/Y sky130_fd_sc_hd__nand2_1
X_4171_ _4175_/A _4171_/B VGND VGND VPWR VPWR _4171_/X sky130_fd_sc_hd__or2_1
X_3122_ _3338_/A _3121_/Y _5080_/Q _5117_/Q VGND VGND VPWR VPWR _3123_/A sky130_fd_sc_hd__o22a_1
XFILLER_67_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3053_ _5072_/Q VGND VGND VPWR VPWR _3330_/A sky130_fd_sc_hd__clkinv_1
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3955_ _3984_/A _3818_/X _3852_/X VGND VGND VPWR VPWR _3956_/A sky130_fd_sc_hd__o21ai_1
X_2906_ _5051_/Q VGND VGND VPWR VPWR _3525_/A sky130_fd_sc_hd__buf_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3886_ _4153_/A VGND VGND VPWR VPWR _3985_/A sky130_fd_sc_hd__clkbuf_2
X_2837_ _2837_/A _2837_/B _2837_/C _2837_/D VGND VGND VPWR VPWR _2840_/B sky130_fd_sc_hd__or4_4
X_2768_ _2768_/A _2821_/B VGND VGND VPWR VPWR _2768_/X sky130_fd_sc_hd__or2_1
X_2699_ _2567_/X _2606_/B _2659_/X VGND VGND VPWR VPWR _2701_/C sky130_fd_sc_hd__o21a_1
X_4507_ _4507_/A _4507_/B VGND VGND VPWR VPWR _4507_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4438_ _4372_/X _4387_/X _4577_/A _4437_/X VGND VGND VPWR VPWR _4546_/A sky130_fd_sc_hd__o31a_2
X_4369_ _4369_/A VGND VGND VPWR VPWR _4632_/B sky130_fd_sc_hd__buf_1
XFILLER_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer50 _3344_/B VGND VGND VPWR VPWR _3404_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3740_ _4601_/A _3740_/B VGND VGND VPWR VPWR _4975_/D sky130_fd_sc_hd__nor2_1
XFILLER_13_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3671_ _3679_/A _3671_/B VGND VGND VPWR VPWR _5005_/D sky130_fd_sc_hd__nor2_1
X_2622_ _2622_/A VGND VGND VPWR VPWR _2777_/A sky130_fd_sc_hd__inv_2
X_2553_ _2560_/A VGND VGND VPWR VPWR _2553_/X sky130_fd_sc_hd__buf_1
X_2484_ _4687_/B _2484_/B VGND VGND VPWR VPWR _2484_/Y sky130_fd_sc_hd__nand2_1
X_4223_ _4250_/A _4084_/X _4118_/X VGND VGND VPWR VPWR _4224_/A sky130_fd_sc_hd__o21ai_1
X_4154_ _4154_/A _4154_/B VGND VGND VPWR VPWR _4155_/C sky130_fd_sc_hd__nand2_1
X_3105_ _5077_/Q _3030_/X _5076_/Q _5113_/Q VGND VGND VPWR VPWR _3105_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4085_ _4981_/Q VGND VGND VPWR VPWR _4086_/B sky130_fd_sc_hd__inv_2
X_3036_ _3036_/A VGND VGND VPWR VPWR _3264_/A sky130_fd_sc_hd__inv_2
XFILLER_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4987_ _5028_/CLK _4987_/D VGND VGND VPWR VPWR _4987_/Q sky130_fd_sc_hd__dfxtp_1
X_3938_ _3938_/A VGND VGND VPWR VPWR _3938_/Y sky130_fd_sc_hd__inv_2
X_3869_ _3602_/B _5036_/Q _3604_/B _5035_/Q VGND VGND VPWR VPWR _3869_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 mdata1 VGND VGND VPWR VPWR _3323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4910_ _5028_/CLK _4910_/D VGND VGND VPWR VPWR _4910_/Q sky130_fd_sc_hd__dfxtp_1
X_4841_ _5028_/CLK _4841_/D VGND VGND VPWR VPWR _4841_/Q sky130_fd_sc_hd__dfxtp_1
X_4772_ _5139_/Q _4772_/D VGND VGND VPWR VPWR _4772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3723_ _3725_/A _3723_/B VGND VGND VPWR VPWR _4982_/D sky130_fd_sc_hd__nor2_1
X_3654_ _3656_/A _3654_/B VGND VGND VPWR VPWR _5013_/D sky130_fd_sc_hd__nor2_1
X_2605_ _2781_/A VGND VGND VPWR VPWR _2606_/B sky130_fd_sc_hd__clkbuf_2
X_3585_ _4932_/Q VGND VGND VPWR VPWR _3586_/B sky130_fd_sc_hd__inv_2
X_2536_ _2543_/A VGND VGND VPWR VPWR _2536_/X sky130_fd_sc_hd__buf_1
X_2467_ _4692_/A _2475_/B _4694_/Y VGND VGND VPWR VPWR _2468_/B sky130_fd_sc_hd__o21ai_1
X_4206_ _4206_/A VGND VGND VPWR VPWR _4206_/Y sky130_fd_sc_hd__inv_2
X_2398_ _4614_/B _2968_/X _4678_/A _2396_/Y _2397_/X VGND VGND VPWR VPWR _2398_/X
+ sky130_fd_sc_hd__o221a_1
X_4137_ _3679_/B _5001_/Q _3683_/B _5000_/Q VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__a211o_1
X_4068_ _3710_/B _4988_/Q _3710_/B _4988_/Q VGND VGND VPWR VPWR _4222_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3019_ _3344_/A _2991_/X _3016_/X _3018_/Y VGND VGND VPWR VPWR _3019_/X sky130_fd_sc_hd__a22o_1
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3370_ _3370_/A VGND VGND VPWR VPWR _4639_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5040_ _5047_/CLK _5040_/D VGND VGND VPWR VPWR _5040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4824_ _4648_/X _4824_/D VGND VGND VPWR VPWR _4824_/Q sky130_fd_sc_hd__dfxtp_1
X_4755_ _2642_/Y _2575_/X _4770_/S VGND VGND VPWR VPWR _4772_/D sky130_fd_sc_hd__mux2_2
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3706_ _3714_/A _3706_/B VGND VGND VPWR VPWR _4990_/D sky130_fd_sc_hd__nor2_1
X_4686_ _4348_/A _3008_/A _4806_/Q _5119_/Q VGND VGND VPWR VPWR _4687_/B sky130_fd_sc_hd__o22a_1
X_3637_ _3645_/A _3637_/B VGND VGND VPWR VPWR _5021_/D sky130_fd_sc_hd__nor2_1
X_3568_ _3568_/A VGND VGND VPWR VPWR _3568_/Y sky130_fd_sc_hd__inv_2
X_2519_ _2519_/A VGND VGND VPWR VPWR _2519_/X sky130_fd_sc_hd__buf_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3499_ input6/X _3498_/X _3494_/Y VGND VGND VPWR VPWR _3500_/A sky130_fd_sc_hd__a21oi_2
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2870_ _2866_/A _3503_/B _3512_/B VGND VGND VPWR VPWR _2870_/Y sky130_fd_sc_hd__a21oi_4
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4540_ _4342_/A _4538_/Y _4339_/A _4538_/A _4539_/X VGND VGND VPWR VPWR _4882_/D
+ sky130_fd_sc_hd__o221a_1
X_4471_ _4823_/Q VGND VGND VPWR VPWR _4605_/B sky130_fd_sc_hd__inv_2
X_3422_ _3422_/A VGND VGND VPWR VPWR _3422_/Y sky130_fd_sc_hd__clkinvlp_2
X_3353_ _3353_/A _3353_/B VGND VGND VPWR VPWR _3354_/B sky130_fd_sc_hd__or2_1
X_3284_ _3057_/A _3283_/Y _3052_/A _3283_/A _3267_/X VGND VGND VPWR VPWR _5110_/D
+ sky130_fd_sc_hd__o221a_1
X_5023_ _5028_/CLK _5023_/D VGND VGND VPWR VPWR _5023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4807_ _2482_/X _4807_/D VGND VGND VPWR VPWR _4807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2999_ _3342_/A _2998_/Y _5084_/Q _5121_/Q VGND VGND VPWR VPWR _3000_/A sky130_fd_sc_hd__o22a_1
X_4738_ _4644_/B _3086_/X _4729_/Y _4643_/B _3100_/Y VGND VGND VPWR VPWR _4738_/X
+ sky130_fd_sc_hd__o32a_1
X_4669_ _4669_/A _4669_/B VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3971_ _3971_/A _3971_/B VGND VGND VPWR VPWR _3971_/Y sky130_fd_sc_hd__nand2_1
X_2922_ _2922_/A _2922_/B _2922_/C VGND VGND VPWR VPWR _2923_/B sky130_fd_sc_hd__nor3_4
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2853_ input4/X _2857_/A VGND VGND VPWR VPWR _3508_/B sky130_fd_sc_hd__or2_2
X_2784_ _2610_/A _2783_/X _2733_/X VGND VGND VPWR VPWR _2785_/D sky130_fd_sc_hd__o21a_1
X_4523_ _4620_/B _4848_/Q _4522_/Y VGND VGND VPWR VPWR _4524_/A sky130_fd_sc_hd__o21ai_1
X_4454_ _4452_/X _4294_/Y _4453_/X VGND VGND VPWR VPWR _4454_/Y sky130_fd_sc_hd__o21ai_1
X_4385_ _4637_/B _4834_/Q _4384_/A _4834_/Q VGND VGND VPWR VPWR _4577_/B sky130_fd_sc_hd__a2bb2o_1
X_3405_ _4176_/A VGND VGND VPWR VPWR _3978_/A sky130_fd_sc_hd__clkbuf_4
X_3336_ _3336_/A _3336_/B VGND VGND VPWR VPWR _3337_/B sky130_fd_sc_hd__or2_1
XFILLER_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5006_ _5047_/CLK _5006_/D VGND VGND VPWR VPWR _5006_/Q sky130_fd_sc_hd__dfxtp_1
X_3267_ _3936_/A VGND VGND VPWR VPWR _3267_/X sky130_fd_sc_hd__buf_2
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3198_ _3212_/A _2985_/B _3134_/Y VGND VGND VPWR VPWR _3199_/B sky130_fd_sc_hd__o21ai_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4170_ _4166_/A _4166_/B _3978_/X _4166_/Y VGND VGND VPWR VPWR _4930_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3121_ _5117_/Q VGND VGND VPWR VPWR _3121_/Y sky130_fd_sc_hd__inv_2
X_3052_ _3052_/A VGND VGND VPWR VPWR _3057_/A sky130_fd_sc_hd__inv_2
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3954_ _3954_/A VGND VGND VPWR VPWR _3958_/A sky130_fd_sc_hd__inv_2
X_3885_ _3748_/Y _3884_/Y _3748_/A _3884_/A _3359_/X VGND VGND VPWR VPWR _4972_/D
+ sky130_fd_sc_hd__o221a_1
X_2905_ _2895_/Y _2897_/A _5050_/Q _2897_/Y _2904_/X VGND VGND VPWR VPWR _2914_/A
+ sky130_fd_sc_hd__a221o_1
X_2836_ _4963_/Q _2777_/A _2778_/A VGND VGND VPWR VPWR _2837_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2767_ _2831_/B VGND VGND VPWR VPWR _2821_/B sky130_fd_sc_hd__buf_1
X_4506_ _4517_/A _4320_/B _4457_/Y VGND VGND VPWR VPWR _4507_/B sky130_fd_sc_hd__o21ai_1
X_2698_ _2698_/A _2698_/B _2698_/C _2698_/D VGND VGND VPWR VPWR _2701_/B sky130_fd_sc_hd__or4_4
X_4437_ _4372_/A _4427_/Y _4372_/X _4433_/X _4436_/X VGND VGND VPWR VPWR _4437_/X
+ sky130_fd_sc_hd__o221a_1
X_4368_ _4800_/Q VGND VGND VPWR VPWR _4369_/A sky130_fd_sc_hd__inv_2
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4299_ _4461_/A _4856_/Q _4461_/A _4856_/Q VGND VGND VPWR VPWR _4488_/A sky130_fd_sc_hd__a2bb2o_1
X_3319_ _3365_/A VGND VGND VPWR VPWR _3319_/X sky130_fd_sc_hd__buf_1
XFILLER_73_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer51 _3334_/B VGND VGND VPWR VPWR _3434_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer40 _3354_/B VGND VGND VPWR VPWR _3374_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3670_ _4894_/Q VGND VGND VPWR VPWR _3671_/B sky130_fd_sc_hd__inv_2
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2621_ _2637_/D _2621_/B _2621_/C _4964_/Q VGND VGND VPWR VPWR _2622_/A sky130_fd_sc_hd__or4b_4
X_2552_ _2547_/A _4728_/B _3318_/C _2548_/A VGND VGND VPWR VPWR _4792_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2483_ _4750_/X _2387_/B _4689_/Y VGND VGND VPWR VPWR _2484_/B sky130_fd_sc_hd__o21ai_1
X_4222_ _4222_/A VGND VGND VPWR VPWR _4226_/A sky130_fd_sc_hd__inv_2
X_4153_ _4153_/A VGND VGND VPWR VPWR _4481_/A sky130_fd_sc_hd__clkbuf_2
X_3104_ _3103_/A _3103_/B _3074_/Y _3077_/X _3103_/X VGND VGND VPWR VPWR _3286_/A
+ sky130_fd_sc_hd__o311a_2
X_4084_ _4084_/A _4084_/B VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__or2_1
X_3035_ _3334_/A _3034_/Y _5076_/Q _5113_/Q VGND VGND VPWR VPWR _3036_/A sky130_fd_sc_hd__o22a_1
XFILLER_55_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4986_ _5028_/CLK _4986_/D VGND VGND VPWR VPWR _4986_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3937_ _3782_/A _3935_/Y _3780_/A _3935_/A _3936_/X VGND VGND VPWR VPWR _4958_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3868_ _4929_/Q _3756_/Y _3867_/X VGND VGND VPWR VPWR _3868_/Y sky130_fd_sc_hd__o21ai_1
X_2819_ _4967_/Q _2783_/X _2798_/X VGND VGND VPWR VPWR _2820_/D sky130_fd_sc_hd__o21a_1
X_3799_ _4915_/Q _3799_/B VGND VGND VPWR VPWR _3799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 reset VGND VGND VPWR VPWR _3370_/A sky130_fd_sc_hd__buf_2
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4840_ _5028_/CLK _4840_/D VGND VGND VPWR VPWR _4840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4771_ _3576_/B _2923_/B _5138_/Q VGND VGND VPWR VPWR _4771_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3722_ _4871_/Q VGND VGND VPWR VPWR _3723_/B sky130_fd_sc_hd__inv_2
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3653_ _4902_/Q VGND VGND VPWR VPWR _3654_/B sky130_fd_sc_hd__inv_2
X_2604_ _2611_/A _2604_/B _2616_/C VGND VGND VPWR VPWR _2781_/A sky130_fd_sc_hd__nor3_4
X_3584_ _3588_/A _3584_/B VGND VGND VPWR VPWR _5044_/D sky130_fd_sc_hd__nor2_1
X_2535_ _2534_/Y _4713_/A _2517_/X _2529_/X VGND VGND VPWR VPWR _4796_/D sky130_fd_sc_hd__o211a_1
X_2466_ _2466_/A VGND VGND VPWR VPWR _2475_/B sky130_fd_sc_hd__inv_2
X_4205_ _4048_/A _4204_/Y _4046_/A _4204_/A _4190_/X VGND VGND VPWR VPWR _4921_/D
+ sky130_fd_sc_hd__o221a_1
X_4136_ _4888_/Q _4036_/Y _4135_/Y VGND VGND VPWR VPWR _4136_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2397_ _4614_/B _2968_/X _4616_/B _2972_/X VGND VGND VPWR VPWR _2397_/X sky130_fd_sc_hd__a211o_1
X_4067_ _4067_/A VGND VGND VPWR VPWR _4069_/A sky130_fd_sc_hd__inv_2
X_3018_ _5085_/Q _2992_/X _3017_/X VGND VGND VPWR VPWR _3018_/Y sky130_fd_sc_hd__o21ai_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4969_ _5018_/CLK _4969_/D VGND VGND VPWR VPWR _4969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4823_ _2410_/X _4823_/D VGND VGND VPWR VPWR _4823_/Q sky130_fd_sc_hd__dfxtp_2
X_4754_ _4754_/A VGND VGND VPWR VPWR _4754_/Y sky130_fd_sc_hd__inv_2
X_3705_ _4879_/Q VGND VGND VPWR VPWR _3706_/B sky130_fd_sc_hd__inv_2
X_4685_ _4807_/Q _5120_/Q _4337_/A _3004_/A VGND VGND VPWR VPWR _4687_/A sky130_fd_sc_hd__o22a_1
X_3636_ _4910_/Q VGND VGND VPWR VPWR _3637_/B sky130_fd_sc_hd__inv_2
X_3567_ _3480_/A _3480_/B _3481_/B _3556_/A VGND VGND VPWR VPWR _5055_/D sky130_fd_sc_hd__a211oi_2
XFILLER_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2518_ _4704_/A _2503_/A _2517_/X _2512_/X VGND VGND VPWR VPWR _4800_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3498_ _3498_/A _3498_/B VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__or2_1
X_2449_ _4616_/B _2972_/X _2448_/Y VGND VGND VPWR VPWR _2451_/B sky130_fd_sc_hd__o21ai_1
XFILLER_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4119_ _3710_/B _4988_/Q _4065_/Y _3708_/B _4989_/Q VGND VGND VPWR VPWR _4119_/X
+ sky130_fd_sc_hd__o32a_1
X_5099_ _3361_/X _5099_/D VGND VGND VPWR VPWR _5099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4470_ _4470_/A VGND VGND VPWR VPWR _4606_/B sky130_fd_sc_hd__clkbuf_2
X_3421_ _3426_/A VGND VGND VPWR VPWR _3421_/X sky130_fd_sc_hd__buf_1
X_3352_ _3352_/A _3352_/B VGND VGND VPWR VPWR _3353_/B sky130_fd_sc_hd__or2_1
X_3283_ _3283_/A VGND VGND VPWR VPWR _3283_/Y sky130_fd_sc_hd__inv_2
X_5022_ _5028_/CLK _5022_/D VGND VGND VPWR VPWR _5022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4806_ _2489_/X _4806_/D VGND VGND VPWR VPWR _4806_/Q sky130_fd_sc_hd__dfxtp_1
X_2998_ _5121_/Q VGND VGND VPWR VPWR _2998_/Y sky130_fd_sc_hd__inv_2
X_4737_ _4737_/A VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__inv_2
X_4668_ _4668_/A _4668_/B VGND VGND VPWR VPWR _4669_/B sky130_fd_sc_hd__nand2_1
X_3619_ _4917_/Q VGND VGND VPWR VPWR _3620_/B sky130_fd_sc_hd__inv_2
X_4599_ _4788_/Q VGND VGND VPWR VPWR _4735_/A sky130_fd_sc_hd__inv_2
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3970_ _3984_/A _3818_/B _3850_/Y VGND VGND VPWR VPWR _3971_/B sky130_fd_sc_hd__o21ai_1
XFILLER_62_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2921_ _5060_/Q _2863_/Y _2868_/X _2874_/Y _2920_/X VGND VGND VPWR VPWR _2922_/B
+ sky130_fd_sc_hd__a2111o_4
XFILLER_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2852_ input2/X input3/X _3503_/B VGND VGND VPWR VPWR _2857_/A sky130_fd_sc_hd__or3_1
X_2783_ _2783_/A VGND VGND VPWR VPWR _2783_/X sky130_fd_sc_hd__clkbuf_2
X_4522_ _4522_/A _4522_/B VGND VGND VPWR VPWR _4522_/Y sky130_fd_sc_hd__nand2_1
X_4453_ _4613_/B _4854_/Q _4452_/X _4294_/Y VGND VGND VPWR VPWR _4453_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3404_ _3404_/A VGND VGND VPWR VPWR _3404_/Y sky130_fd_sc_hd__inv_2
X_4384_ _4384_/A VGND VGND VPWR VPWR _4637_/B sky130_fd_sc_hd__buf_1
X_3335_ _3335_/A _3335_/B VGND VGND VPWR VPWR _3336_/B sky130_fd_sc_hd__or2_1
X_3266_ _3266_/A VGND VGND VPWR VPWR _3266_/Y sky130_fd_sc_hd__inv_2
X_5005_ _5047_/CLK _5005_/D VGND VGND VPWR VPWR _5005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3197_ _3197_/A VGND VGND VPWR VPWR _3197_/X sky130_fd_sc_hd__buf_1
XFILLER_53_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3120_ _5080_/Q VGND VGND VPWR VPWR _3338_/A sky130_fd_sc_hd__clkinv_1
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3051_ _3331_/A _3049_/Y _5073_/Q _3050_/X VGND VGND VPWR VPWR _3052_/A sky130_fd_sc_hd__o22a_1
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ _3952_/Y _3859_/A _3939_/X _3948_/X VGND VGND VPWR VPWR _4953_/D sky130_fd_sc_hd__o211a_1
X_3884_ _3884_/A VGND VGND VPWR VPWR _3884_/Y sky130_fd_sc_hd__inv_2
X_2904_ _2899_/X input8/X _2902_/Y _2902_/A _2903_/Y VGND VGND VPWR VPWR _2904_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_31_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2835_ _2756_/A _2774_/A _2775_/A VGND VGND VPWR VPWR _2837_/C sky130_fd_sc_hd__o21a_1
X_2766_ _2766_/A _2766_/B _2766_/C _2766_/D VGND VGND VPWR VPWR _2766_/X sky130_fd_sc_hd__or4_4
X_4505_ _4505_/A VGND VGND VPWR VPWR _4507_/A sky130_fd_sc_hd__inv_2
X_2697_ _2736_/A _2624_/B _2590_/D VGND VGND VPWR VPWR _2698_/D sky130_fd_sc_hd__o21a_1
X_4436_ _4630_/B _4840_/Q _4357_/Y _4629_/B _4841_/Q VGND VGND VPWR VPWR _4436_/X
+ sky130_fd_sc_hd__o32a_1
X_4367_ _4367_/A VGND VGND VPWR VPWR _4371_/A sky130_fd_sc_hd__inv_2
X_3318_ _3316_/X _3318_/B _3318_/C VGND VGND VPWR VPWR _5102_/D sky130_fd_sc_hd__and3b_1
XFILLER_58_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4298_ _4818_/Q VGND VGND VPWR VPWR _4461_/A sky130_fd_sc_hd__inv_2
X_3249_ _3269_/A VGND VGND VPWR VPWR _3249_/X sky130_fd_sc_hd__buf_1
XFILLER_66_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer30 _3339_/B VGND VGND VPWR VPWR _3420_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer41 _3328_/B VGND VGND VPWR VPWR _3451_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer52 _3342_/B VGND VGND VPWR VPWR _3411_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2620_ _4951_/Q _2632_/B _2620_/C _2620_/D VGND VGND VPWR VPWR _2637_/D sky130_fd_sc_hd__or4_4
X_2551_ _2560_/A VGND VGND VPWR VPWR _2551_/X sky130_fd_sc_hd__buf_1
X_2482_ _2497_/A VGND VGND VPWR VPWR _2482_/X sky130_fd_sc_hd__buf_1
X_4221_ _4219_/Y _4125_/A _4220_/X _4215_/X VGND VGND VPWR VPWR _4916_/D sky130_fd_sc_hd__o211a_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4152_ _4014_/Y _4150_/Y _4014_/A _4150_/A _4151_/X VGND VGND VPWR VPWR _4935_/D
+ sky130_fd_sc_hd__o221a_1
X_3103_ _3103_/A _3103_/B _3103_/C _3290_/A VGND VGND VPWR VPWR _3103_/X sky130_fd_sc_hd__or4_4
XFILLER_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4083_ _4083_/A _4250_/B VGND VGND VPWR VPWR _4084_/B sky130_fd_sc_hd__or2_1
X_3034_ _5113_/Q VGND VGND VPWR VPWR _3034_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4985_ _5028_/CLK _4985_/D VGND VGND VPWR VPWR _4985_/Q sky130_fd_sc_hd__dfxtp_1
X_3936_ _3936_/A VGND VGND VPWR VPWR _3936_/X sky130_fd_sc_hd__clkbuf_2
X_3867_ _3595_/B _5039_/Q _4929_/Q _3756_/Y VGND VGND VPWR VPWR _3867_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2818_ _4970_/Q _2781_/X _2796_/X VGND VGND VPWR VPWR _2820_/C sky130_fd_sc_hd__o21a_1
X_3798_ _5026_/Q VGND VGND VPWR VPWR _3799_/B sky130_fd_sc_hd__inv_2
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2749_ _4944_/Q _2726_/X _2707_/X VGND VGND VPWR VPWR _2752_/B sky130_fd_sc_hd__o21a_1
X_4419_ _4419_/A VGND VGND VPWR VPWR _4592_/A sky130_fd_sc_hd__inv_2
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4770_ _2840_/X _2831_/X _4770_/S VGND VGND VPWR VPWR _4787_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3721_ _3725_/A _3721_/B VGND VGND VPWR VPWR _4983_/D sky130_fd_sc_hd__nor2_1
X_3652_ _3656_/A _3652_/B VGND VGND VPWR VPWR _5014_/D sky130_fd_sc_hd__nor2_1
X_3583_ _4933_/Q VGND VGND VPWR VPWR _3584_/B sky130_fd_sc_hd__inv_2
X_2603_ _4961_/Q _2610_/A _2621_/B _2603_/D VGND VGND VPWR VPWR _2616_/C sky130_fd_sc_hd__or4_4
X_2534_ _4741_/X VGND VGND VPWR VPWR _2534_/Y sky130_fd_sc_hd__inv_2
X_2465_ _4750_/X _2391_/A _4692_/B VGND VGND VPWR VPWR _2466_/A sky130_fd_sc_hd__o21ai_1
X_4204_ _4204_/A VGND VGND VPWR VPWR _4204_/Y sky130_fd_sc_hd__inv_2
X_2396_ _4312_/X _2977_/X _2395_/X VGND VGND VPWR VPWR _2396_/Y sky130_fd_sc_hd__o21ai_2
X_4135_ _3685_/B _4999_/Q _3687_/B _4998_/Q VGND VGND VPWR VPWR _4135_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4066_ _4878_/Q _4065_/B _4065_/Y VGND VGND VPWR VPWR _4067_/A sky130_fd_sc_hd__a21oi_2
X_3017_ _5085_/Q _2992_/X _5084_/Q _5121_/Q VGND VGND VPWR VPWR _3017_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4968_ _5018_/CLK _4968_/D VGND VGND VPWR VPWR _4968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3919_ _3923_/A _3923_/B VGND VGND VPWR VPWR _3924_/B sky130_fd_sc_hd__or2_1
X_4899_ _5047_/CLK _4899_/D VGND VGND VPWR VPWR _4899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4822_ _2415_/X _4822_/D VGND VGND VPWR VPWR _4822_/Q sky130_fd_sc_hd__dfxtp_1
X_4753_ _4628_/B _3121_/Y _4804_/Q _5117_/Q VGND VGND VPWR VPWR _4754_/A sky130_fd_sc_hd__o22a_1
X_3704_ _3726_/A VGND VGND VPWR VPWR _3714_/A sky130_fd_sc_hd__clkbuf_2
X_4684_ _4684_/A _4684_/B VGND VGND VPWR VPWR _4692_/A sky130_fd_sc_hd__or2_1
X_3635_ _3669_/A VGND VGND VPWR VPWR _3645_/A sky130_fd_sc_hd__clkbuf_2
X_3566_ _3481_/A _3481_/B _3482_/A _3559_/X VGND VGND VPWR VPWR _5056_/D sky130_fd_sc_hd__o211a_1
X_3497_ _2880_/Y _3496_/A _5063_/Q _3496_/Y VGND VGND VPWR VPWR _3551_/A sky130_fd_sc_hd__o22a_1
X_2517_ _3165_/A VGND VGND VPWR VPWR _2517_/X sky130_fd_sc_hd__clkbuf_2
X_2448_ _4672_/B _2448_/B VGND VGND VPWR VPWR _2448_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4118_ _3717_/B _4985_/Q _4084_/A _4116_/Y _4117_/X VGND VGND VPWR VPWR _4118_/X
+ sky130_fd_sc_hd__o221a_1
X_5098_ _3365_/X _5098_/D VGND VGND VPWR VPWR _5098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4049_ _3699_/B _4993_/Q _3699_/B _4993_/Q VGND VGND VPWR VPWR _4050_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3420_ _3339_/A _3420_/A2 _3401_/X _3417_/Y VGND VGND VPWR VPWR _5081_/D sky130_fd_sc_hd__a211oi_1
X_3351_ _3351_/A _3351_/B VGND VGND VPWR VPWR _3352_/B sky130_fd_sc_hd__or2_1
X_3282_ _3330_/A _3054_/Y _3281_/X VGND VGND VPWR VPWR _3283_/A sky130_fd_sc_hd__o21ai_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5021_ _5028_/CLK _5021_/D VGND VGND VPWR VPWR _5021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4805_ _2491_/X _4805_/D VGND VGND VPWR VPWR _4805_/Q sky130_fd_sc_hd__dfxtp_1
X_2997_ _5084_/Q VGND VGND VPWR VPWR _3342_/A sky130_fd_sc_hd__clkinv_1
X_4736_ _4645_/B _3091_/Y _4735_/X VGND VGND VPWR VPWR _4737_/A sky130_fd_sc_hd__o21ai_2
X_4667_ _4819_/Q _5132_/Q _4666_/Y VGND VGND VPWR VPWR _4668_/B sky130_fd_sc_hd__a21oi_2
X_3618_ _3622_/A _3618_/B VGND VGND VPWR VPWR _5029_/D sky130_fd_sc_hd__nor2_1
X_4598_ _4788_/Q _4414_/Y _4416_/X _3165_/X _4417_/Y VGND VGND VPWR VPWR _4864_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3549_ _5061_/Q _3546_/Y _3548_/X VGND VGND VPWR VPWR _3549_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2920_ _3487_/A _2876_/X _2919_/Y VGND VGND VPWR VPWR _2920_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2851_ _3501_/A _3502_/B VGND VGND VPWR VPWR _3503_/B sky130_fd_sc_hd__or2_4
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2782_ _4967_/Q _2781_/X _2731_/X VGND VGND VPWR VPWR _2785_/C sky130_fd_sc_hd__o21a_1
Xclkbuf_0_mclk1 mclk1 VGND VGND VPWR VPWR clkbuf_0_mclk1/X sky130_fd_sc_hd__clkbuf_16
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4521_ _4450_/C _4528_/B _4353_/Y VGND VGND VPWR VPWR _4522_/B sky130_fd_sc_hd__o21ai_1
X_4452_ _4817_/Q VGND VGND VPWR VPWR _4452_/X sky130_fd_sc_hd__clkbuf_2
X_3403_ _3413_/A VGND VGND VPWR VPWR _3403_/X sky130_fd_sc_hd__buf_1
X_4383_ _4796_/Q VGND VGND VPWR VPWR _4384_/A sky130_fd_sc_hd__inv_2
X_3334_ _3334_/A _3334_/B VGND VGND VPWR VPWR _3335_/B sky130_fd_sc_hd__or2_1
X_3265_ _3334_/A _3034_/Y _3264_/X VGND VGND VPWR VPWR _3266_/A sky130_fd_sc_hd__o21ai_1
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_mclk1 clkbuf_0_mclk1/X VGND VGND VPWR VPWR _5139_/CLK sky130_fd_sc_hd__clkbuf_1
X_5004_ _5047_/CLK _5004_/D VGND VGND VPWR VPWR _5004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3196_ _2951_/A _3178_/A _3186_/X _3189_/X VGND VGND VPWR VPWR _5129_/D sky130_fd_sc_hd__o211a_1
XFILLER_26_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4719_ _4401_/A _3064_/A _4794_/Q _5107_/Q VGND VGND VPWR VPWR _4720_/A sky130_fd_sc_hd__o22a_1
XFILLER_1_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3050_ _5110_/Q VGND VGND VPWR VPWR _3050_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3952_ _3952_/A VGND VGND VPWR VPWR _3952_/Y sky130_fd_sc_hd__inv_2
X_3883_ _3582_/B _5045_/Q _3888_/B VGND VGND VPWR VPWR _3884_/A sky130_fd_sc_hd__o21ai_1
X_2903_ _2903_/A input8/X VGND VGND VPWR VPWR _2903_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2834_ _4951_/Q _2791_/X _2772_/A VGND VGND VPWR VPWR _2837_/B sky130_fd_sc_hd__o21a_1
X_2765_ _4963_/Q _2718_/X _2733_/X VGND VGND VPWR VPWR _2766_/D sky130_fd_sc_hd__o21a_1
X_4504_ _4503_/Y _4490_/A _4264_/X _4497_/X VGND VGND VPWR VPWR _4891_/D sky130_fd_sc_hd__o211a_1
X_2696_ _4943_/Q _2630_/B _2590_/C VGND VGND VPWR VPWR _2698_/C sky130_fd_sc_hd__o21a_1
X_4435_ _4803_/Q VGND VGND VPWR VPWR _4629_/B sky130_fd_sc_hd__inv_2
X_4366_ _4631_/B _4839_/Q _4364_/X _4365_/Y VGND VGND VPWR VPWR _4367_/A sky130_fd_sc_hd__o22a_1
X_3317_ _4500_/A VGND VGND VPWR VPWR _3318_/C sky130_fd_sc_hd__clkbuf_2
X_4297_ _4503_/A _4297_/B VGND VGND VPWR VPWR _4305_/A sky130_fd_sc_hd__or2_1
X_3248_ _3368_/A VGND VGND VPWR VPWR _3269_/A sky130_fd_sc_hd__buf_1
XFILLER_39_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer20 _3343_/B VGND VGND VPWR VPWR _3412_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_3179_ _2965_/A _3189_/B _3132_/Y VGND VGND VPWR VPWR _3180_/B sky130_fd_sc_hd__o21ai_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer31 _3331_/B VGND VGND VPWR VPWR _3447_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer42 _3340_/B VGND VGND VPWR VPWR _3417_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer53 _3356_/B VGND VGND VPWR VPWR _3366_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2550_ _4722_/Y _2548_/Y _4728_/A _3165_/X _2549_/Y VGND VGND VPWR VPWR _4793_/D
+ sky130_fd_sc_hd__o311a_1
X_2481_ _4683_/A _2466_/A _2450_/X _2475_/X VGND VGND VPWR VPWR _4808_/D sky130_fd_sc_hd__o211a_1
X_4220_ _4562_/A VGND VGND VPWR VPWR _4220_/X sky130_fd_sc_hd__clkbuf_2
X_4151_ _4269_/A VGND VGND VPWR VPWR _4151_/X sky130_fd_sc_hd__clkbuf_2
X_3102_ _3083_/Y _3308_/B _3308_/A _3101_/X VGND VGND VPWR VPWR _3290_/A sky130_fd_sc_hd__o31a_1
X_4082_ _3723_/B _4982_/Q _3723_/B _4982_/Q VGND VGND VPWR VPWR _4250_/B sky130_fd_sc_hd__a2bb2o_1
X_3033_ _5076_/Q VGND VGND VPWR VPWR _3334_/A sky130_fd_sc_hd__clkinv_1
XFILLER_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4984_ _5028_/CLK _4984_/D VGND VGND VPWR VPWR _4984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3935_ _3935_/A VGND VGND VPWR VPWR _3935_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3866_ _3777_/Y _3797_/X _3952_/A _3865_/X VGND VGND VPWR VPWR _3923_/A sky130_fd_sc_hd__o22a_2
X_2817_ _2817_/A _2817_/B _2817_/C _2817_/D VGND VGND VPWR VPWR _2820_/B sky130_fd_sc_hd__or4_4
X_3797_ _3606_/B _5034_/Q _3609_/B _5033_/Q _3796_/X VGND VGND VPWR VPWR _3797_/X
+ sky130_fd_sc_hd__o221a_1
X_2748_ _2703_/A _2705_/X _2693_/X VGND VGND VPWR VPWR _2752_/A sky130_fd_sc_hd__o21a_1
X_2679_ _2679_/A _2679_/B _2679_/C _2679_/D VGND VGND VPWR VPWR _2679_/X sky130_fd_sc_hd__or4_1
X_4418_ _4645_/B _4827_/Q _4417_/Y VGND VGND VPWR VPWR _4419_/A sky130_fd_sc_hd__o21ai_2
X_4349_ _4624_/B _4845_/Q _4625_/B _4844_/Q VGND VGND VPWR VPWR _4349_/X sky130_fd_sc_hd__a211o_1
XFILLER_27_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3720_ _4872_/Q VGND VGND VPWR VPWR _3721_/B sky130_fd_sc_hd__inv_2
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3651_ _4903_/Q VGND VGND VPWR VPWR _3652_/B sky130_fd_sc_hd__inv_2
X_3582_ _3588_/A _3582_/B VGND VGND VPWR VPWR _5045_/D sky130_fd_sc_hd__nor2_1
X_2602_ _4962_/Q _4963_/Q VGND VGND VPWR VPWR _2621_/B sky130_fd_sc_hd__or2_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2533_ _2543_/A VGND VGND VPWR VPWR _2533_/X sky130_fd_sc_hd__buf_1
X_2464_ _2474_/A VGND VGND VPWR VPWR _2464_/X sky130_fd_sc_hd__buf_1
XFILLER_68_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4203_ _3697_/B _4994_/Q _4202_/X VGND VGND VPWR VPWR _4204_/A sky130_fd_sc_hd__o21ai_1
X_2395_ _4312_/X _2977_/X _4812_/Q _5125_/Q VGND VGND VPWR VPWR _2395_/X sky130_fd_sc_hd__a22o_1
X_4134_ _4892_/Q _4022_/Y _4133_/X VGND VGND VPWR VPWR _4134_/Y sky130_fd_sc_hd__o21ai_1
X_4065_ _4878_/Q _4065_/B VGND VGND VPWR VPWR _4065_/Y sky130_fd_sc_hd__nor2_1
X_3016_ _3129_/C _3016_/B VGND VGND VPWR VPWR _3016_/X sky130_fd_sc_hd__or2_1
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4967_ _5018_/CLK _4967_/D VGND VGND VPWR VPWR _4967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3918_ _3913_/A _3913_/B _3462_/X _3913_/Y VGND VGND VPWR VPWR _4963_/D sky130_fd_sc_hd__o211a_1
X_4898_ _5047_/CLK _4898_/D VGND VGND VPWR VPWR _4898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3849_ _3639_/B _5020_/Q _3641_/B _5019_/Q VGND VGND VPWR VPWR _3849_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_59_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4821_ _2419_/X _4821_/D VGND VGND VPWR VPWR _4821_/Q sky130_fd_sc_hd__dfxtp_2
X_4752_ _4752_/A VGND VGND VPWR VPWR _4752_/Y sky130_fd_sc_hd__inv_2
X_4683_ _4683_/A VGND VGND VPWR VPWR _4684_/B sky130_fd_sc_hd__inv_2
X_3703_ _3703_/A _3703_/B VGND VGND VPWR VPWR _4991_/D sky130_fd_sc_hd__nor2_1
X_3634_ _3634_/A _3634_/B VGND VGND VPWR VPWR _5022_/D sky130_fd_sc_hd__nor2_1
X_3565_ _3483_/A _3483_/B _3484_/B _3559_/X VGND VGND VPWR VPWR _5057_/D sky130_fd_sc_hd__o211a_1
X_2516_ _2519_/A VGND VGND VPWR VPWR _2516_/X sky130_fd_sc_hd__buf_1
X_3496_ _3496_/A VGND VGND VPWR VPWR _3496_/Y sky130_fd_sc_hd__inv_2
X_2447_ _2462_/A _4678_/B _2396_/Y VGND VGND VPWR VPWR _2448_/B sky130_fd_sc_hd__o21ai_1
XFILLER_68_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4117_ _3717_/B _4985_/Q _3719_/B _4984_/Q VGND VGND VPWR VPWR _4117_/X sky130_fd_sc_hd__a211o_1
X_5097_ _3369_/X _5097_/D VGND VGND VPWR VPWR _5097_/Q sky130_fd_sc_hd__dfxtp_1
X_4048_ _4048_/A _4206_/A VGND VGND VPWR VPWR _4131_/C sky130_fd_sc_hd__or2_1
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3350_ _3350_/A _3350_/B VGND VGND VPWR VPWR _3351_/B sky130_fd_sc_hd__or2_1
X_3281_ _3286_/A _3281_/B VGND VGND VPWR VPWR _3281_/X sky130_fd_sc_hd__or2_1
X_5020_ _5028_/CLK _5020_/D VGND VGND VPWR VPWR _5020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4804_ _2497_/X _4804_/D VGND VGND VPWR VPWR _4804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2996_ _2996_/A VGND VGND VPWR VPWR _3001_/A sky130_fd_sc_hd__inv_2
X_4735_ _4735_/A _4735_/B _4735_/C VGND VGND VPWR VPWR _4735_/X sky130_fd_sc_hd__or3_1
X_4666_ _4819_/Q _5132_/Q VGND VGND VPWR VPWR _4666_/Y sky130_fd_sc_hd__nor2_1
X_3617_ _4918_/Q VGND VGND VPWR VPWR _3618_/B sky130_fd_sc_hd__inv_2
X_4597_ _4419_/A _4596_/Y _4562_/X _4592_/X VGND VGND VPWR VPWR _4865_/D sky130_fd_sc_hd__o211a_1
X_3548_ _5058_/Q _3547_/Y _5058_/Q _3547_/Y VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3479_ _3479_/A _3568_/A VGND VGND VPWR VPWR _3480_/B sky130_fd_sc_hd__or2_2
XFILLER_69_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2850_ _2850_/A _3518_/B VGND VGND VPWR VPWR _3502_/B sky130_fd_sc_hd__or2_2
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _2781_/A VGND VGND VPWR VPWR _2781_/X sky130_fd_sc_hd__clkbuf_2
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4520_ _4520_/A VGND VGND VPWR VPWR _4528_/B sky130_fd_sc_hd__inv_2
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4451_ _4322_/Y _4355_/X _4546_/A _4450_/X VGND VGND VPWR VPWR _4517_/A sky130_fd_sc_hd__o22a_2
X_3402_ _3345_/A _3402_/A2 _3401_/X _3397_/Y VGND VGND VPWR VPWR _5087_/D sky130_fd_sc_hd__a211oi_2
X_4382_ _4382_/A VGND VGND VPWR VPWR _4386_/A sky130_fd_sc_hd__inv_2
X_3333_ _3333_/A _3333_/B VGND VGND VPWR VPWR _3334_/B sky130_fd_sc_hd__or2_1
X_3264_ _3264_/A _3264_/B VGND VGND VPWR VPWR _3264_/X sky130_fd_sc_hd__or2_1
X_5003_ _5047_/CLK _5003_/D VGND VGND VPWR VPWR _5003_/Q sky130_fd_sc_hd__dfxtp_1
X_3195_ _3197_/A VGND VGND VPWR VPWR _3195_/X sky130_fd_sc_hd__buf_1
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2979_ _2979_/A VGND VGND VPWR VPWR _2984_/A sky130_fd_sc_hd__inv_2
X_4718_ _4718_/A VGND VGND VPWR VPWR _4740_/A sky130_fd_sc_hd__inv_2
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4649_ _4824_/Q _5137_/Q _4604_/B _2930_/Y VGND VGND VPWR VPWR _4649_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3951_ _3860_/A _3950_/Y _3857_/A _3950_/A _3936_/X VGND VGND VPWR VPWR _4954_/D
+ sky130_fd_sc_hd__o221a_1
X_2902_ _2902_/A VGND VGND VPWR VPWR _2902_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3882_ _3887_/A _3887_/B VGND VGND VPWR VPWR _3888_/B sky130_fd_sc_hd__or2_1
XFILLER_31_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2833_ _4957_/Q _2770_/A _2758_/A VGND VGND VPWR VPWR _2837_/A sky130_fd_sc_hd__o21a_1
X_2764_ _4966_/Q _2716_/X _2731_/X VGND VGND VPWR VPWR _2766_/C sky130_fd_sc_hd__o21a_1
X_4503_ _4503_/A VGND VGND VPWR VPWR _4503_/Y sky130_fd_sc_hd__inv_2
X_2695_ _4940_/Q _2651_/X _2590_/B VGND VGND VPWR VPWR _2698_/B sky130_fd_sc_hd__o21a_1
X_4434_ _4434_/A VGND VGND VPWR VPWR _4630_/B sky130_fd_sc_hd__clkbuf_2
X_4365_ _4839_/Q VGND VGND VPWR VPWR _4365_/Y sky130_fd_sc_hd__inv_2
X_3316_ _3324_/A _3096_/B _3096_/C VGND VGND VPWR VPWR _3316_/X sky130_fd_sc_hd__o21a_1
X_4296_ _4296_/A VGND VGND VPWR VPWR _4297_/B sky130_fd_sc_hd__inv_2
X_3247_ _3384_/A VGND VGND VPWR VPWR _3368_/A sky130_fd_sc_hd__buf_1
XFILLER_73_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer21 _3343_/B VGND VGND VPWR VPWR _3409_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer10 _3327_/B VGND VGND VPWR VPWR _3454_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_3178_ _3178_/A VGND VGND VPWR VPWR _3189_/B sky130_fd_sc_hd__inv_2
XFILLER_54_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer43 _3330_/B VGND VGND VPWR VPWR _3446_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer32 _3331_/B VGND VGND VPWR VPWR _3443_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer54 _3326_/B VGND VGND VPWR VPWR rebuffer1/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2480_ _2497_/A VGND VGND VPWR VPWR _2480_/X sky130_fd_sc_hd__buf_1
X_4150_ _4150_/A VGND VGND VPWR VPWR _4150_/Y sky130_fd_sc_hd__inv_2
X_3101_ _3324_/D _3086_/X _3081_/Y _3325_/A _3100_/Y VGND VGND VPWR VPWR _3101_/X
+ sky130_fd_sc_hd__o32a_1
X_4081_ _4081_/A VGND VGND VPWR VPWR _4083_/A sky130_fd_sc_hd__inv_2
X_3032_ _3032_/A VGND VGND VPWR VPWR _3037_/A sky130_fd_sc_hd__inv_2
XFILLER_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4983_ _5028_/CLK _4983_/D VGND VGND VPWR VPWR _4983_/Q sky130_fd_sc_hd__dfxtp_1
X_3934_ _3614_/B _5031_/Q _3933_/X VGND VGND VPWR VPWR _3935_/A sky130_fd_sc_hd__o21ai_1
X_3865_ _3865_/A _3865_/B _3865_/C _3928_/A VGND VGND VPWR VPWR _3865_/X sky130_fd_sc_hd__or4b_4
X_2816_ _2567_/X _2777_/X _2778_/X VGND VGND VPWR VPWR _2817_/D sky130_fd_sc_hd__o21a_1
X_3796_ _3609_/B _5033_/Q _3793_/X _3795_/Y VGND VGND VPWR VPWR _3796_/X sky130_fd_sc_hd__a22o_1
X_2747_ _2821_/A _2722_/X _2723_/X VGND VGND VPWR VPWR _2755_/A sky130_fd_sc_hd__o21a_1
X_2678_ _2786_/A _2613_/B _2663_/X VGND VGND VPWR VPWR _2679_/D sky130_fd_sc_hd__o21a_1
X_4417_ _4788_/Q _4414_/Y _4416_/X VGND VGND VPWR VPWR _4417_/Y sky130_fd_sc_hd__o21ai_1
X_4348_ _4348_/A VGND VGND VPWR VPWR _4625_/B sky130_fd_sc_hd__clkbuf_2
X_4279_ _4823_/Q _4279_/B VGND VGND VPWR VPWR _4279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3650_ _3656_/A _3825_/A VGND VGND VPWR VPWR _5015_/D sky130_fd_sc_hd__nor2_1
X_3581_ _4934_/Q VGND VGND VPWR VPWR _3582_/B sky130_fd_sc_hd__inv_2
X_2601_ _4964_/Q VGND VGND VPWR VPWR _2610_/A sky130_fd_sc_hd__clkbuf_2
Xrebuffer1 rebuffer1/A VGND VGND VPWR VPWR _3463_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_2532_ _4714_/A _2531_/Y _4711_/A _2531_/A _2495_/X VGND VGND VPWR VPWR _4797_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4202_ _4206_/A _4202_/B VGND VGND VPWR VPWR _4202_/X sky130_fd_sc_hd__or2_1
X_2463_ _2462_/Y _4676_/A _2450_/X _2457_/X VGND VGND VPWR VPWR _4812_/D sky130_fd_sc_hd__o211a_1
X_2394_ _4452_/X _2952_/X _2393_/X VGND VGND VPWR VPWR _2394_/Y sky130_fd_sc_hd__o21ai_1
X_4133_ _3677_/B _5002_/Q _4892_/Q _4022_/Y VGND VGND VPWR VPWR _4133_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4064_ _4989_/Q VGND VGND VPWR VPWR _4065_/B sky130_fd_sc_hd__inv_2
X_3015_ _3341_/A _3004_/X _3125_/A _3013_/Y _3014_/X VGND VGND VPWR VPWR _3016_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4966_ _5018_/CLK _4966_/D VGND VGND VPWR VPWR _4966_/Q sky130_fd_sc_hd__dfxtp_1
X_3917_ _3916_/A _3915_/Y _3916_/Y _3915_/A _3902_/X VGND VGND VPWR VPWR _4964_/D
+ sky130_fd_sc_hd__o221a_1
X_4897_ _5047_/CLK _4897_/D VGND VGND VPWR VPWR _4897_/Q sky130_fd_sc_hd__dfxtp_1
X_3848_ _4913_/Q _3804_/Y _3847_/Y VGND VGND VPWR VPWR _3848_/Y sky130_fd_sc_hd__o21ai_1
X_3779_ _4921_/Q _3778_/Y _3611_/B _5032_/Q VGND VGND VPWR VPWR _3780_/A sky130_fd_sc_hd__o22a_1
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4820_ _2425_/X _4820_/D VGND VGND VPWR VPWR _4820_/Q sky130_fd_sc_hd__dfxtp_1
X_4751_ _4343_/X _3011_/X _4626_/B _3117_/Y VGND VGND VPWR VPWR _4752_/A sky130_fd_sc_hd__o22a_1
XFILLER_14_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4682_ _4333_/A _2998_/Y _4808_/Q _5121_/Q VGND VGND VPWR VPWR _4683_/A sky130_fd_sc_hd__o22a_1
X_3702_ _4880_/Q VGND VGND VPWR VPWR _3703_/B sky130_fd_sc_hd__inv_2
X_3633_ _4911_/Q VGND VGND VPWR VPWR _3634_/B sky130_fd_sc_hd__inv_2
X_3564_ _3484_/A _3484_/B _3562_/Y _3556_/A VGND VGND VPWR VPWR _5058_/D sky130_fd_sc_hd__a211oi_1
X_2515_ _4705_/A _2514_/Y _4702_/A _2514_/A _2495_/X VGND VGND VPWR VPWR _4801_/D
+ sky130_fd_sc_hd__o221a_1
X_3495_ _3490_/Y _3494_/Y _3498_/A _2859_/A VGND VGND VPWR VPWR _3496_/A sky130_fd_sc_hd__o22a_1
X_2446_ _2453_/A VGND VGND VPWR VPWR _2446_/X sky130_fd_sc_hd__buf_1
X_4116_ _4872_/Q _4079_/Y _4115_/Y VGND VGND VPWR VPWR _4116_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5096_ _3373_/X _5096_/D VGND VGND VPWR VPWR _5096_/Q sky130_fd_sc_hd__dfxtp_1
X_4047_ _3697_/B _4994_/Q _3697_/B _4994_/Q VGND VGND VPWR VPWR _4206_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4949_ _5018_/CLK _4949_/D VGND VGND VPWR VPWR _4949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3280_ _3289_/A VGND VGND VPWR VPWR _3280_/X sky130_fd_sc_hd__buf_1
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4803_ _2501_/X _4803_/D VGND VGND VPWR VPWR _4803_/Q sky130_fd_sc_hd__dfxtp_2
X_2995_ _5085_/Q _2992_/X _3343_/A _2994_/Y VGND VGND VPWR VPWR _2996_/A sky130_fd_sc_hd__o22a_1
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4734_ _4789_/Q _5102_/Q _4645_/B _3091_/Y VGND VGND VPWR VPWR _4735_/C sky130_fd_sc_hd__a22o_1
X_4665_ _4818_/Q _5131_/Q _4461_/A _2960_/A VGND VGND VPWR VPWR _4668_/A sky130_fd_sc_hd__o22a_1
X_4596_ _4596_/A VGND VGND VPWR VPWR _4596_/Y sky130_fd_sc_hd__inv_2
X_3616_ _3622_/A _3616_/B VGND VGND VPWR VPWR _5030_/D sky130_fd_sc_hd__nor2_1
X_3547_ _2866_/A _3503_/X _3513_/Y VGND VGND VPWR VPWR _3547_/Y sky130_fd_sc_hd__a21oi_1
X_3478_ _3478_/A _3478_/B VGND VGND VPWR VPWR _3568_/A sky130_fd_sc_hd__or2_1
XFILLER_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2429_ _2462_/A _4678_/X _2398_/X VGND VGND VPWR VPWR _2430_/A sky130_fd_sc_hd__o21ai_1
XFILLER_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5079_ _3424_/X _5079_/D VGND VGND VPWR VPWR _5079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ _2780_/A _2780_/B _2780_/C _2780_/D VGND VGND VPWR VPWR _2785_/B sky130_fd_sc_hd__or4_4
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ _4450_/A _4450_/B _4450_/C _4522_/A VGND VGND VPWR VPWR _4450_/X sky130_fd_sc_hd__or4b_4
X_3401_ _4639_/A VGND VGND VPWR VPWR _3401_/X sky130_fd_sc_hd__buf_2
X_4381_ _4636_/B _4835_/Q _4379_/X _4380_/Y VGND VGND VPWR VPWR _4382_/A sky130_fd_sc_hd__o22a_1
X_3332_ _3332_/A _3332_/B VGND VGND VPWR VPWR _3333_/B sky130_fd_sc_hd__or2_1
X_3263_ _3269_/A VGND VGND VPWR VPWR _3263_/X sky130_fd_sc_hd__buf_1
X_5002_ _5047_/CLK _5002_/D VGND VGND VPWR VPWR _5002_/Q sky130_fd_sc_hd__dfxtp_1
X_3194_ _2957_/B _3191_/Y _2956_/A _3191_/A _3193_/X VGND VGND VPWR VPWR _5130_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2978_ _3347_/A _2976_/Y _5089_/Q _2977_/X VGND VGND VPWR VPWR _2979_/A sky130_fd_sc_hd__o22a_1
X_4717_ _4795_/Q _5108_/Q _4716_/Y VGND VGND VPWR VPWR _4718_/A sky130_fd_sc_hd__a21oi_2
X_4648_ _4648_/A VGND VGND VPWR VPWR _4648_/X sky130_fd_sc_hd__buf_1
X_4579_ _4579_/A VGND VGND VPWR VPWR _4582_/A sky130_fd_sc_hd__inv_2
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3950_ _3950_/A VGND VGND VPWR VPWR _3950_/Y sky130_fd_sc_hd__inv_2
X_2901_ _2900_/Y input9/X _2900_/Y input9/X VGND VGND VPWR VPWR _2902_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3881_ _3744_/Y _3880_/A _3744_/A _3880_/Y _3359_/X VGND VGND VPWR VPWR _4973_/D
+ sky130_fd_sc_hd__o221a_1
X_2832_ _4966_/Q _2787_/X _2788_/X VGND VGND VPWR VPWR _2840_/A sky130_fd_sc_hd__o21a_1
XFILLER_31_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2763_ _2763_/A _2763_/B _2763_/C _2763_/D VGND VGND VPWR VPWR _2766_/B sky130_fd_sc_hd__or4_4
X_4502_ _4297_/B _4499_/Y _4296_/A _4499_/A _4501_/X VGND VGND VPWR VPWR _4892_/D
+ sky130_fd_sc_hd__o221a_1
X_2694_ _2643_/A _2638_/X _2693_/X VGND VGND VPWR VPWR _2698_/A sky130_fd_sc_hd__o21a_1
X_4433_ _4634_/B _4837_/Q _4387_/A _4430_/Y _4432_/X VGND VGND VPWR VPWR _4433_/X
+ sky130_fd_sc_hd__o221a_1
X_4364_ _4801_/Q VGND VGND VPWR VPWR _4364_/X sky130_fd_sc_hd__clkbuf_2
X_4295_ _4612_/B _4855_/Q _4817_/Q _4294_/Y VGND VGND VPWR VPWR _4296_/A sky130_fd_sc_hd__o22a_1
X_3315_ _3365_/A VGND VGND VPWR VPWR _3315_/X sky130_fd_sc_hd__buf_1
X_3246_ _3246_/A VGND VGND VPWR VPWR _3384_/A sky130_fd_sc_hd__buf_1
XFILLER_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer11 _3327_/B VGND VGND VPWR VPWR _3457_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3177_ _3212_/A _2985_/X _3136_/X VGND VGND VPWR VPWR _3178_/A sky130_fd_sc_hd__o21ai_1
Xrebuffer22 _3345_/B VGND VGND VPWR VPWR _3407_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer55 _3326_/B VGND VGND VPWR VPWR rebuffer2/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer33 _3336_/B VGND VGND VPWR VPWR _3427_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer44 _3323_/A VGND VGND VPWR VPWR _3471_/B2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3100_ _5104_/Q VGND VGND VPWR VPWR _3100_/Y sky130_fd_sc_hd__inv_2
X_4080_ _3721_/B _4983_/Q _4872_/Q _4079_/Y VGND VGND VPWR VPWR _4081_/A sky130_fd_sc_hd__o22a_1
X_3031_ _3335_/A _3029_/Y _5077_/Q _3030_/X VGND VGND VPWR VPWR _3032_/A sky130_fd_sc_hd__o22a_1
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4982_ _5028_/CLK _4982_/D VGND VGND VPWR VPWR _4982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3933_ _3938_/A _3933_/B VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__or2_1
X_3864_ _3609_/B _5033_/Q _3608_/A _5033_/Q VGND VGND VPWR VPWR _3928_/A sky130_fd_sc_hd__o2bb2a_1
X_2815_ _2736_/A _2774_/X _2775_/X VGND VGND VPWR VPWR _2817_/C sky130_fd_sc_hd__o21a_1
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3795_ _4921_/Q _3778_/Y _3794_/Y VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__o21ai_1
X_2746_ _2746_/A _2756_/B VGND VGND VPWR VPWR _2746_/X sky130_fd_sc_hd__or2_1
XFILLER_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2677_ _4956_/Q VGND VGND VPWR VPWR _2786_/A sky130_fd_sc_hd__clkbuf_2
X_4416_ _4645_/B _4827_/Q _4789_/Q _4415_/Y VGND VGND VPWR VPWR _4416_/X sky130_fd_sc_hd__o22a_1
X_4347_ _4343_/X _4344_/Y _4346_/X VGND VGND VPWR VPWR _4347_/Y sky130_fd_sc_hd__o21ai_1
X_4278_ _4861_/Q VGND VGND VPWR VPWR _4279_/B sky130_fd_sc_hd__inv_2
X_3229_ _3229_/A VGND VGND VPWR VPWR _3229_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2600_ _4968_/Q _4970_/Q _2600_/C VGND VGND VPWR VPWR _2604_/B sky130_fd_sc_hd__or3_4
X_3580_ _3588_/A _3580_/B VGND VGND VPWR VPWR _5046_/D sky130_fd_sc_hd__nor2_1
Xrebuffer2 rebuffer2/A VGND VGND VPWR VPWR _3456_/A sky130_fd_sc_hd__dlygate4sd1_1
X_2531_ _2531_/A VGND VGND VPWR VPWR _2531_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2462_ _2462_/A VGND VGND VPWR VPWR _2462_/Y sky130_fd_sc_hd__inv_2
X_4201_ _4197_/A _4197_/B _4177_/X _4197_/Y VGND VGND VPWR VPWR _4922_/D sky130_fd_sc_hd__o211a_1
X_2393_ _4816_/Q _5129_/Q _4452_/X _2952_/X VGND VGND VPWR VPWR _2393_/X sky130_fd_sc_hd__a22o_1
X_4132_ _4043_/Y _4063_/X _4219_/A _4131_/X VGND VGND VPWR VPWR _4192_/A sky130_fd_sc_hd__o22a_2
XFILLER_68_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4063_ _3689_/B _4997_/Q _3692_/B _4996_/Q _4062_/X VGND VGND VPWR VPWR _4063_/X
+ sky130_fd_sc_hd__o221a_1
X_3014_ _3341_/A _3004_/X _3340_/A _3008_/X VGND VGND VPWR VPWR _3014_/X sky130_fd_sc_hd__a211o_1
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4965_ _5018_/CLK _4965_/D VGND VGND VPWR VPWR _4965_/Q sky130_fd_sc_hd__dfxtp_1
X_3916_ _3916_/A VGND VGND VPWR VPWR _3916_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4896_ _5047_/CLK _4896_/D VGND VGND VPWR VPWR _4896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ _3630_/B _5024_/Q _3632_/B _5023_/Q VGND VGND VPWR VPWR _3847_/Y sky130_fd_sc_hd__o22ai_1
X_3778_ _5032_/Q VGND VGND VPWR VPWR _3778_/Y sky130_fd_sc_hd__inv_2
X_2729_ _2756_/A _2712_/X _2713_/X VGND VGND VPWR VPWR _2730_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4750_ _4706_/X _4715_/X _4741_/X _4749_/X VGND VGND VPWR VPWR _4750_/X sky130_fd_sc_hd__o31a_2
X_4681_ _4681_/A VGND VGND VPWR VPWR _4684_/A sky130_fd_sc_hd__inv_2
X_3701_ _3703_/A _3701_/B VGND VGND VPWR VPWR _4992_/D sky130_fd_sc_hd__nor2_1
X_3632_ _3634_/A _3632_/B VGND VGND VPWR VPWR _5023_/D sky130_fd_sc_hd__nor2_1
X_3563_ _5059_/Q _3562_/Y _3486_/B _3559_/X VGND VGND VPWR VPWR _5059_/D sky130_fd_sc_hd__o211a_1
X_2514_ _2514_/A VGND VGND VPWR VPWR _2514_/Y sky130_fd_sc_hd__inv_2
X_3494_ _3498_/A _3494_/B VGND VGND VPWR VPWR _3494_/Y sky130_fd_sc_hd__nor2_1
X_2445_ _4661_/A _2430_/A _2417_/X _2440_/X VGND VGND VPWR VPWR _4816_/D sky130_fd_sc_hd__o211a_1
XFILLER_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4115_ _3721_/B _4983_/Q _3723_/B _4982_/Q VGND VGND VPWR VPWR _4115_/Y sky130_fd_sc_hd__o22ai_1
X_5095_ _3377_/X _5095_/D VGND VGND VPWR VPWR _5095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4046_ _4046_/A VGND VGND VPWR VPWR _4048_/A sky130_fd_sc_hd__inv_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4948_ _5018_/CLK _4948_/D VGND VGND VPWR VPWR _4948_/Q sky130_fd_sc_hd__dfxtp_1
X_4879_ _5028_/CLK _4879_/D VGND VGND VPWR VPWR _4879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4802_ _2509_/X _4802_/D VGND VGND VPWR VPWR _4802_/Q sky130_fd_sc_hd__dfxtp_1
X_2994_ _5122_/Q VGND VGND VPWR VPWR _2994_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4733_ _4733_/A VGND VGND VPWR VPWR _4733_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4664_ _4664_/A _4664_/B VGND VGND VPWR VPWR _4669_/A sky130_fd_sc_hd__or2_1
X_4595_ _4410_/Y _4594_/Y _4410_/A _4594_/A _4575_/X VGND VGND VPWR VPWR _4866_/D
+ sky130_fd_sc_hd__o221a_1
X_3615_ _4919_/Q VGND VGND VPWR VPWR _3616_/B sky130_fd_sc_hd__inv_2
X_3546_ input5/X _3508_/X _3498_/X VGND VGND VPWR VPWR _3546_/Y sky130_fd_sc_hd__a21boi_1
X_3477_ _5052_/Q _3477_/B VGND VGND VPWR VPWR _3478_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2428_ _2428_/A VGND VGND VPWR VPWR _2428_/X sky130_fd_sc_hd__buf_1
XFILLER_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5078_ _3426_/X _5078_/D VGND VGND VPWR VPWR _5078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4029_ _4894_/Q _4028_/B _4028_/Y VGND VGND VPWR VPWR _4030_/A sky130_fd_sc_hd__a21oi_2
XFILLER_71_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3400_ _3413_/A VGND VGND VPWR VPWR _3400_/X sky130_fd_sc_hd__buf_1
X_4380_ _4835_/Q VGND VGND VPWR VPWR _4380_/Y sky130_fd_sc_hd__inv_2
X_3331_ _3331_/A _3331_/B VGND VGND VPWR VPWR _3332_/B sky130_fd_sc_hd__or2_1
X_3262_ _3256_/A _3256_/B _3258_/X _3256_/Y VGND VGND VPWR VPWR _5115_/D sky130_fd_sc_hd__o211a_1
X_5001_ _5047_/CLK _5001_/D VGND VGND VPWR VPWR _5001_/Q sky130_fd_sc_hd__dfxtp_1
X_3193_ _3936_/A VGND VGND VPWR VPWR _3193_/X sky130_fd_sc_hd__buf_2
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2977_ _5126_/Q VGND VGND VPWR VPWR _2977_/X sky130_fd_sc_hd__clkbuf_2
X_4716_ _4795_/Q _5108_/Q VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__nor2_1
X_4647_ _4647_/A _4647_/B VGND VGND VPWR VPWR _4825_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4578_ _4578_/A _4578_/B _4578_/C VGND VGND VPWR VPWR _4871_/D sky130_fd_sc_hd__and3_1
X_3529_ input9/X _3522_/B _3523_/B VGND VGND VPWR VPWR _3529_/X sky130_fd_sc_hd__a21bo_1
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2900_ _5049_/Q VGND VGND VPWR VPWR _2900_/Y sky130_fd_sc_hd__inv_2
X_3880_ _3880_/A VGND VGND VPWR VPWR _3880_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2831_ _2831_/A _2831_/B VGND VGND VPWR VPWR _2831_/X sky130_fd_sc_hd__or2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2762_ _2801_/A _2712_/X _2713_/X VGND VGND VPWR VPWR _2763_/D sky130_fd_sc_hd__o21a_1
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4501_ _4575_/A VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__buf_2
XANTENNA_0 dec_rate[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2693_ _2758_/A VGND VGND VPWR VPWR _2693_/X sky130_fd_sc_hd__buf_1
X_4432_ _4634_/B _4837_/Q _4635_/B _4836_/Q VGND VGND VPWR VPWR _4432_/X sky130_fd_sc_hd__a211o_1
XFILLER_6_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4363_ _4801_/Q VGND VGND VPWR VPWR _4631_/B sky130_fd_sc_hd__inv_2
X_4294_ _4855_/Q VGND VGND VPWR VPWR _4294_/Y sky130_fd_sc_hd__inv_2
X_3314_ _3368_/A VGND VGND VPWR VPWR _3365_/A sky130_fd_sc_hd__buf_1
X_3245_ _3124_/A _3244_/Y _3119_/A _3244_/A _3193_/X VGND VGND VPWR VPWR _5118_/D
+ sky130_fd_sc_hd__o221a_1
Xrebuffer12 _3357_/B VGND VGND VPWR VPWR _3367_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_3176_ _3197_/A VGND VGND VPWR VPWR _3176_/X sky130_fd_sc_hd__buf_1
XFILLER_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer45 _3332_/B VGND VGND VPWR VPWR _3440_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer34 _3335_/B VGND VGND VPWR VPWR _3436_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer23 _3345_/B VGND VGND VPWR VPWR _3402_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3030_ _5114_/Q VGND VGND VPWR VPWR _3030_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ _5018_/CLK _4981_/D VGND VGND VPWR VPWR _4981_/Q sky130_fd_sc_hd__dfxtp_1
X_3932_ _3928_/A _3928_/B _3462_/X _3928_/Y VGND VGND VPWR VPWR _4959_/D sky130_fd_sc_hd__o211a_1
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3863_ _3863_/A VGND VGND VPWR VPWR _3865_/B sky130_fd_sc_hd__inv_2
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2814_ _2691_/A _2791_/X _2772_/X VGND VGND VPWR VPWR _2817_/B sky130_fd_sc_hd__o21a_1
X_3794_ _3611_/B _5032_/Q _3614_/B _5031_/Q VGND VGND VPWR VPWR _3794_/Y sky130_fd_sc_hd__o22ai_1
X_2745_ _2745_/A _2745_/B _2745_/C _2745_/D VGND VGND VPWR VPWR _2745_/X sky130_fd_sc_hd__or4_4
X_2676_ _2821_/A _2606_/B _2659_/X VGND VGND VPWR VPWR _2679_/C sky130_fd_sc_hd__o21a_1
X_4415_ _4827_/Q VGND VGND VPWR VPWR _4415_/Y sky130_fd_sc_hd__inv_2
X_4346_ _4805_/Q _4344_/Y _4804_/Q _4345_/Y VGND VGND VPWR VPWR _4346_/X sky130_fd_sc_hd__a22o_1
X_4277_ _4277_/A VGND VGND VPWR VPWR _4277_/Y sky130_fd_sc_hd__inv_2
X_3228_ _3342_/A _2998_/Y _3227_/X VGND VGND VPWR VPWR _3229_/A sky130_fd_sc_hd__o21ai_1
XFILLER_27_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3159_ _3356_/A _2937_/X _3158_/X VGND VGND VPWR VPWR _3160_/A sky130_fd_sc_hd__o21ai_1
XFILLER_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer3 _3324_/B VGND VGND VPWR VPWR _3471_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_2530_ _4637_/B _3054_/Y _2529_/X VGND VGND VPWR VPWR _2531_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2461_ _2474_/A VGND VGND VPWR VPWR _2461_/X sky130_fd_sc_hd__buf_1
X_4200_ _4131_/B _4199_/Y _4129_/A _4199_/A _4190_/X VGND VGND VPWR VPWR _4923_/D
+ sky130_fd_sc_hd__o221a_1
X_2392_ _4679_/Y _4696_/X _4750_/X _2391_/X VGND VGND VPWR VPWR _2462_/A sky130_fd_sc_hd__o22a_2
XFILLER_68_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4131_ _4131_/A _4131_/B _4131_/C _4197_/A VGND VGND VPWR VPWR _4131_/X sky130_fd_sc_hd__or4b_4
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4062_ _3692_/B _4996_/Q _4059_/X _4061_/Y VGND VGND VPWR VPWR _4062_/X sky130_fd_sc_hd__a22o_1
X_3013_ _5081_/Q _3011_/X _3012_/X VGND VGND VPWR VPWR _3013_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4964_ _5018_/CLK _4964_/D VGND VGND VPWR VPWR _4964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3915_ _3915_/A VGND VGND VPWR VPWR _3915_/Y sky130_fd_sc_hd__inv_2
X_4895_ _5047_/CLK _4895_/D VGND VGND VPWR VPWR _4895_/Q sky130_fd_sc_hd__dfxtp_1
X_3846_ _3845_/A _3986_/A _3827_/Y _3828_/X _3845_/X VGND VGND VPWR VPWR _3984_/A
+ sky130_fd_sc_hd__o311a_2
X_3777_ _4923_/Q _3777_/B VGND VGND VPWR VPWR _3777_/Y sky130_fd_sc_hd__nor2_1
X_2728_ _2636_/B _2709_/X _2710_/X VGND VGND VPWR VPWR _2730_/C sky130_fd_sc_hd__o21a_1
X_2659_ _2796_/A VGND VGND VPWR VPWR _2659_/X sky130_fd_sc_hd__buf_1
X_4329_ _4809_/Q VGND VGND VPWR VPWR _4622_/B sky130_fd_sc_hd__inv_2
XFILLER_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3700_ _4881_/Q VGND VGND VPWR VPWR _3701_/B sky130_fd_sc_hd__inv_2
X_4680_ _4327_/X _5122_/Q _4622_/B _2994_/Y VGND VGND VPWR VPWR _4681_/A sky130_fd_sc_hd__o22a_1
X_3631_ _4912_/Q VGND VGND VPWR VPWR _3632_/B sky130_fd_sc_hd__inv_2
X_3562_ _3562_/A VGND VGND VPWR VPWR _3562_/Y sky130_fd_sc_hd__inv_2
X_2513_ _4632_/B _3034_/Y _2512_/X VGND VGND VPWR VPWR _2514_/A sky130_fd_sc_hd__o21ai_1
XFILLER_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3493_ _3508_/A VGND VGND VPWR VPWR _3498_/A sky130_fd_sc_hd__clkbuf_2
X_2444_ _2453_/A VGND VGND VPWR VPWR _2444_/X sky130_fd_sc_hd__buf_1
X_4114_ _4876_/Q _4070_/Y _4113_/Y VGND VGND VPWR VPWR _4114_/Y sky130_fd_sc_hd__o21ai_1
X_5094_ _3379_/X _5094_/D VGND VGND VPWR VPWR _5094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4045_ _4884_/Q _4044_/Y _3695_/B _4995_/Q VGND VGND VPWR VPWR _4046_/A sky130_fd_sc_hd__o22a_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4947_ _5018_/CLK _4947_/D VGND VGND VPWR VPWR _4947_/Q sky130_fd_sc_hd__dfxtp_1
X_4878_ _5028_/CLK _4878_/D VGND VGND VPWR VPWR _4878_/Q sky130_fd_sc_hd__dfxtp_1
X_3829_ _3824_/A _5016_/Q _3824_/Y VGND VGND VPWR VPWR _3831_/A sky130_fd_sc_hd__a21oi_2
XFILLER_79_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2993_ _5085_/Q VGND VGND VPWR VPWR _3343_/A sky130_fd_sc_hd__clkinv_1
X_4801_ _2511_/X _4801_/D VGND VGND VPWR VPWR _4801_/Q sky130_fd_sc_hd__dfxtp_1
X_4732_ _4420_/A _3086_/A _4790_/Q _5103_/Q VGND VGND VPWR VPWR _4733_/A sky130_fd_sc_hd__o22a_1
X_4663_ _4663_/A VGND VGND VPWR VPWR _4664_/B sky130_fd_sc_hd__inv_2
X_3614_ _3622_/A _3614_/B VGND VGND VPWR VPWR _5031_/D sky130_fd_sc_hd__nor2_1
X_4594_ _4594_/A VGND VGND VPWR VPWR _4594_/Y sky130_fd_sc_hd__inv_2
X_3545_ _5062_/Q _3500_/A _3488_/A _3500_/Y _3544_/X VGND VGND VPWR VPWR _3551_/B
+ sky130_fd_sc_hd__a221o_1
X_3476_ _3476_/A VGND VGND VPWR VPWR _3477_/B sky130_fd_sc_hd__inv_2
X_2427_ _2426_/Y _4659_/A _2417_/X _2420_/X VGND VGND VPWR VPWR _4820_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5077_ _3430_/X _5077_/D VGND VGND VPWR VPWR _5077_/Q sky130_fd_sc_hd__dfxtp_1
X_4028_ _4894_/Q _4028_/B VGND VGND VPWR VPWR _4028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3330_ _3330_/A _3330_/B VGND VGND VPWR VPWR _3331_/B sky130_fd_sc_hd__or2_1
X_5000_ _5047_/CLK _5000_/D VGND VGND VPWR VPWR _5000_/Q sky130_fd_sc_hd__dfxtp_1
X_3261_ _3269_/A VGND VGND VPWR VPWR _3261_/X sky130_fd_sc_hd__buf_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3192_ _4500_/A VGND VGND VPWR VPWR _3936_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2976_ _5126_/Q VGND VGND VPWR VPWR _2976_/Y sky130_fd_sc_hd__inv_2
X_4715_ _4715_/A _4715_/B VGND VGND VPWR VPWR _4715_/X sky130_fd_sc_hd__or2_1
X_4646_ _4647_/A _4735_/A VGND VGND VPWR VPWR _4826_/D sky130_fd_sc_hd__nor2_1
X_4577_ _4577_/A _4577_/B VGND VGND VPWR VPWR _4578_/C sky130_fd_sc_hd__nand2_1
XFILLER_1_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3528_ _5049_/Q _3527_/Y _5049_/Q _3527_/Y VGND VGND VPWR VPWR _3531_/B sky130_fd_sc_hd__o2bb2a_1
X_3459_ _3459_/A VGND VGND VPWR VPWR _4648_/A sky130_fd_sc_hd__buf_1
XFILLER_69_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5129_ _3195_/X _5129_/D VGND VGND VPWR VPWR _5129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2830_ _2830_/A _2830_/B _2830_/C _2830_/D VGND VGND VPWR VPWR _2830_/X sky130_fd_sc_hd__or4_1
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2761_ _2680_/A _2709_/X _2710_/X VGND VGND VPWR VPWR _2763_/C sky130_fd_sc_hd__o21a_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2692_ _2768_/A _2645_/X _2647_/X VGND VGND VPWR VPWR _2701_/A sky130_fd_sc_hd__o21a_1
X_4500_ _4500_/A VGND VGND VPWR VPWR _4575_/A sky130_fd_sc_hd__buf_1
XANTENNA_1 dec_rate[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4431_ _4431_/A VGND VGND VPWR VPWR _4635_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4362_ _4362_/A _4548_/A VGND VGND VPWR VPWR _4372_/A sky130_fd_sc_hd__or2_1
X_4293_ _4817_/Q VGND VGND VPWR VPWR _4612_/B sky130_fd_sc_hd__inv_2
X_3313_ _3098_/A _3088_/A _3287_/X _3308_/X VGND VGND VPWR VPWR _5103_/D sky130_fd_sc_hd__o211a_1
X_3244_ _3244_/A VGND VGND VPWR VPWR _3244_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3175_ _3225_/A VGND VGND VPWR VPWR _3197_/A sky130_fd_sc_hd__buf_1
Xrebuffer24 _3329_/B VGND VGND VPWR VPWR _3452_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer35 _3335_/B VGND VGND VPWR VPWR _3432_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer46 _3337_/B VGND VGND VPWR VPWR _3428_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer13 _3357_/B VGND VGND VPWR VPWR _3364_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2959_ _5131_/Q VGND VGND VPWR VPWR _2960_/A sky130_fd_sc_hd__inv_2
X_4629_ _4632_/A _4629_/B VGND VGND VPWR VPWR _4841_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4980_ _5018_/CLK _4980_/D VGND VGND VPWR VPWR _4980_/Q sky130_fd_sc_hd__dfxtp_1
X_3931_ _3865_/B _3930_/Y _3863_/A _3930_/A _3902_/X VGND VGND VPWR VPWR _4960_/D
+ sky130_fd_sc_hd__o221a_1
X_3862_ _4923_/Q _3777_/B _3777_/Y VGND VGND VPWR VPWR _3863_/A sky130_fd_sc_hd__a21oi_2
X_2813_ _2768_/A _2770_/X _2758_/X VGND VGND VPWR VPWR _2817_/A sky130_fd_sc_hd__o21a_1
X_3793_ _3865_/C _3793_/B VGND VGND VPWR VPWR _3793_/X sky130_fd_sc_hd__or2_1
X_2744_ _2567_/X _2718_/X _2733_/X VGND VGND VPWR VPWR _2745_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2675_ _4959_/Q VGND VGND VPWR VPWR _2821_/A sky130_fd_sc_hd__clkbuf_2
X_4414_ _4826_/Q VGND VGND VPWR VPWR _4414_/Y sky130_fd_sc_hd__inv_2
X_4345_ _4842_/Q VGND VGND VPWR VPWR _4345_/Y sky130_fd_sc_hd__inv_2
X_4276_ _4824_/Q _4862_/Q _4824_/Q _4862_/Q VGND VGND VPWR VPWR _4277_/A sky130_fd_sc_hd__a2bb2o_1
X_3227_ _3227_/A _3227_/B VGND VGND VPWR VPWR _3227_/X sky130_fd_sc_hd__or2_1
X_3158_ _3163_/A _3158_/B VGND VGND VPWR VPWR _3158_/X sky130_fd_sc_hd__or2_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3089_ _5065_/Q VGND VGND VPWR VPWR _3324_/C sky130_fd_sc_hd__clkinvlp_2
XFILLER_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer4 _3324_/B VGND VGND VPWR VPWR _3469_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_2460_ _4677_/A _2459_/Y _4674_/A _2459_/A _2423_/X VGND VGND VPWR VPWR _4813_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2391_ _2391_/A _2391_/B _4692_/A _2468_/A VGND VGND VPWR VPWR _2391_/X sky130_fd_sc_hd__or4b_4
X_4130_ _3692_/B _4996_/Q _3691_/A _4996_/Q VGND VGND VPWR VPWR _4197_/A sky130_fd_sc_hd__o2bb2a_1
X_4061_ _4884_/Q _4044_/Y _4060_/Y VGND VGND VPWR VPWR _4061_/Y sky130_fd_sc_hd__o21ai_1
X_3012_ _5081_/Q _3011_/X _5080_/Q _5117_/Q VGND VGND VPWR VPWR _3012_/X sky130_fd_sc_hd__a22o_1
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4963_ _5018_/CLK _4963_/D VGND VGND VPWR VPWR _4963_/Q sky130_fd_sc_hd__dfxtp_1
X_3914_ _3599_/B _5037_/Q _3913_/Y VGND VGND VPWR VPWR _3915_/A sky130_fd_sc_hd__o21ai_1
X_4894_ _5047_/CLK _4894_/D VGND VGND VPWR VPWR _4894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3845_ _3845_/A _3986_/A _3845_/C _3987_/A VGND VGND VPWR VPWR _3845_/X sky130_fd_sc_hd__or4_4
X_3776_ _5034_/Q VGND VGND VPWR VPWR _3777_/B sky130_fd_sc_hd__inv_2
X_2727_ _4942_/Q _2726_/X _2707_/X VGND VGND VPWR VPWR _2730_/B sky130_fd_sc_hd__o21a_1
X_2658_ _2658_/A VGND VGND VPWR VPWR _2796_/A sky130_fd_sc_hd__inv_2
XFILLER_59_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2589_ _2778_/A VGND VGND VPWR VPWR _2590_/D sky130_fd_sc_hd__buf_1
X_4328_ _4847_/Q VGND VGND VPWR VPWR _4328_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4259_ _4255_/A _4255_/B _4220_/X _4255_/Y VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__o211a_1
XFILLER_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3630_ _3634_/A _3630_/B VGND VGND VPWR VPWR _5024_/D sky130_fd_sc_hd__nor2_1
X_3561_ _3486_/A _3486_/B _3558_/Y _3576_/B VGND VGND VPWR VPWR _5060_/D sky130_fd_sc_hd__a211oi_1
X_2512_ _4705_/B _2512_/B VGND VGND VPWR VPWR _2512_/X sky130_fd_sc_hd__or2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3492_ _3518_/A VGND VGND VPWR VPWR _3508_/A sky130_fd_sc_hd__buf_1
X_2443_ _4664_/B _2442_/Y _4663_/A _2442_/A _2423_/X VGND VGND VPWR VPWR _4817_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4113_ _3712_/B _4987_/Q _3714_/B _4986_/Q VGND VGND VPWR VPWR _4113_/Y sky130_fd_sc_hd__o22ai_1
X_5093_ _3382_/X _5093_/D VGND VGND VPWR VPWR _5093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4044_ _4995_/Q VGND VGND VPWR VPWR _4044_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4946_ _5018_/CLK _4946_/D VGND VGND VPWR VPWR _4946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4877_ _5028_/CLK _4877_/D VGND VGND VPWR VPWR _4877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3828_ _3645_/B _5017_/Q _3820_/Y _3643_/B _5018_/Q VGND VGND VPWR VPWR _3828_/X
+ sky130_fd_sc_hd__o32a_1
X_3759_ _3909_/A _3759_/B VGND VGND VPWR VPWR _3766_/A sky130_fd_sc_hd__or2_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4800_ _2516_/X _4800_/D VGND VGND VPWR VPWR _4800_/Q sky130_fd_sc_hd__dfxtp_1
X_2992_ _5122_/Q VGND VGND VPWR VPWR _2992_/X sky130_fd_sc_hd__clkbuf_2
X_4731_ _4731_/A VGND VGND VPWR VPWR _4731_/Y sky130_fd_sc_hd__inv_2
X_4662_ _4452_/X _5130_/Q _4612_/B _2954_/Y VGND VGND VPWR VPWR _4663_/A sky130_fd_sc_hd__o22a_1
X_3613_ _4920_/Q VGND VGND VPWR VPWR _3614_/B sky130_fd_sc_hd__inv_2
X_4593_ _4644_/B _4828_/Q _4592_/X VGND VGND VPWR VPWR _4594_/A sky130_fd_sc_hd__o21ai_1
X_3544_ _3544_/A _3544_/B _3544_/C VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__or3_1
X_3475_ _5051_/Q _3574_/A VGND VGND VPWR VPWR _3476_/A sky130_fd_sc_hd__nand2_1
X_2426_ _2426_/A VGND VGND VPWR VPWR _2426_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5076_ _3433_/X _5076_/D VGND VGND VPWR VPWR _5076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4027_ _5005_/Q VGND VGND VPWR VPWR _4028_/B sky130_fd_sc_hd__inv_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4929_ _5047_/CLK _4929_/D VGND VGND VPWR VPWR _4929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3260_ _3259_/A _3259_/B _3258_/X _3259_/Y VGND VGND VPWR VPWR _5116_/D sky130_fd_sc_hd__o211a_1
X_3191_ _3191_/A VGND VGND VPWR VPWR _3191_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4714_ _4714_/A _4714_/B VGND VGND VPWR VPWR _4715_/B sky130_fd_sc_hd__or2_1
X_2975_ _5089_/Q VGND VGND VPWR VPWR _3347_/A sky130_fd_sc_hd__clkinv_1
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4645_ _4647_/A _4645_/B VGND VGND VPWR VPWR _4827_/D sky130_fd_sc_hd__nor2_1
X_4576_ _4386_/A _4574_/Y _4382_/A _4574_/A _4575_/X VGND VGND VPWR VPWR _4872_/D
+ sky130_fd_sc_hd__o221a_1
X_3527_ _2899_/X input8/X _2903_/Y VGND VGND VPWR VPWR _3527_/Y sky130_fd_sc_hd__o21ai_1
X_3458_ _3458_/A VGND VGND VPWR VPWR _3459_/A sky130_fd_sc_hd__buf_1
XFILLER_39_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3389_ _3396_/A VGND VGND VPWR VPWR _3389_/X sky130_fd_sc_hd__buf_1
X_2409_ _3459_/A VGND VGND VPWR VPWR _2428_/A sky130_fd_sc_hd__buf_1
X_5128_ _3197_/X _5128_/D VGND VGND VPWR VPWR _5128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5059_ _5063_/CLK _5059_/D VGND VGND VPWR VPWR _5059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2760_ _2636_/B _2726_/X _2707_/X VGND VGND VPWR VPWR _2763_/B sky130_fd_sc_hd__o21a_1
X_2691_ _2691_/A _2691_/B VGND VGND VPWR VPWR _2691_/X sky130_fd_sc_hd__or2_1
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4430_ _4379_/X _4380_/Y _4429_/Y VGND VGND VPWR VPWR _4430_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_2 _4827_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4361_ _4434_/A _4840_/Q _4434_/A _4840_/Q VGND VGND VPWR VPWR _4548_/A sky130_fd_sc_hd__a2bb2o_1
X_4292_ _4613_/B _4854_/Q _4291_/A _4854_/Q VGND VGND VPWR VPWR _4503_/A sky130_fd_sc_hd__a2bb2o_1
X_3312_ _3312_/A VGND VGND VPWR VPWR _3312_/X sky130_fd_sc_hd__buf_1
X_3243_ _3338_/A _3121_/Y _3242_/X VGND VGND VPWR VPWR _3244_/A sky130_fd_sc_hd__o21ai_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3174_ _3173_/Y _2947_/A _3165_/X _3168_/X VGND VGND VPWR VPWR _5133_/D sky130_fd_sc_hd__o211a_1
Xrebuffer25 _3329_/B VGND VGND VPWR VPWR _3449_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer36 _3338_/B VGND VGND VPWR VPWR _3422_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer14 _3349_/B VGND VGND VPWR VPWR _3393_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer47 _3337_/B VGND VGND VPWR VPWR _3425_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2958_ _5094_/Q VGND VGND VPWR VPWR _3352_/A sky130_fd_sc_hd__clkinvlp_4
X_2889_ _2889_/A VGND VGND VPWR VPWR _2889_/Y sky130_fd_sc_hd__inv_2
X_4628_ _4632_/A _4628_/B VGND VGND VPWR VPWR _4842_/D sky130_fd_sc_hd__nor2_1
X_4559_ _4559_/A VGND VGND VPWR VPWR _4559_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3930_ _3930_/A VGND VGND VPWR VPWR _3930_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3861_ _3861_/A _3861_/B VGND VGND VPWR VPWR _3865_/A sky130_fd_sc_hd__or2_1
X_2812_ _2610_/A _2787_/X _2788_/X VGND VGND VPWR VPWR _2820_/A sky130_fd_sc_hd__o21a_1
X_3792_ _3616_/B _5030_/Q _3861_/A _3790_/Y _3791_/X VGND VGND VPWR VPWR _3793_/B
+ sky130_fd_sc_hd__o221a_1
X_2743_ _2610_/A _2716_/X _2731_/X VGND VGND VPWR VPWR _2745_/C sky130_fd_sc_hd__o21a_1
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2674_ _2674_/A _2674_/B _2674_/C _2674_/D VGND VGND VPWR VPWR _2679_/B sky130_fd_sc_hd__or4_4
X_4413_ _4789_/Q VGND VGND VPWR VPWR _4645_/B sky130_fd_sc_hd__inv_2
X_4344_ _4843_/Q VGND VGND VPWR VPWR _4344_/Y sky130_fd_sc_hd__inv_2
X_4275_ _4601_/A _4275_/B VGND VGND VPWR VPWR _4900_/D sky130_fd_sc_hd__nor2_1
X_3226_ _3241_/A VGND VGND VPWR VPWR _3226_/X sky130_fd_sc_hd__buf_1
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3157_ _3172_/A VGND VGND VPWR VPWR _3157_/X sky130_fd_sc_hd__buf_1
XFILLER_54_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3088_ _3088_/A VGND VGND VPWR VPWR _3308_/B sky130_fd_sc_hd__inv_2
XFILLER_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer5 _3324_/B VGND VGND VPWR VPWR _3468_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_2390_ _4810_/Q _5123_/Q _4326_/A _2991_/A VGND VGND VPWR VPWR _2468_/A sky130_fd_sc_hd__o22a_1
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4060_ _3695_/B _4995_/Q _3697_/B _4994_/Q VGND VGND VPWR VPWR _4060_/Y sky130_fd_sc_hd__o22ai_1
X_3011_ _5118_/Q VGND VGND VPWR VPWR _3011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4962_ _5018_/CLK _4962_/D VGND VGND VPWR VPWR _4962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4893_ _5047_/CLK _4893_/D VGND VGND VPWR VPWR _4893_/Q sky130_fd_sc_hd__dfxtp_1
X_3913_ _3913_/A _3913_/B VGND VGND VPWR VPWR _3913_/Y sky130_fd_sc_hd__nand2_1
X_3844_ _3835_/Y _4004_/A _4000_/A _3843_/X VGND VGND VPWR VPWR _3987_/A sky130_fd_sc_hd__o31a_1
X_3775_ _3775_/A _3775_/B VGND VGND VPWR VPWR _3775_/X sky130_fd_sc_hd__or2_1
X_2726_ _2791_/A VGND VGND VPWR VPWR _2726_/X sky130_fd_sc_hd__clkbuf_2
X_2657_ _4958_/Q VGND VGND VPWR VPWR _2811_/A sky130_fd_sc_hd__clkbuf_2
X_2588_ _2588_/A VGND VGND VPWR VPWR _2778_/A sky130_fd_sc_hd__inv_2
X_4327_ _4809_/Q VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4258_ _4111_/A _4257_/Y _4088_/A _4257_/A _4229_/X VGND VGND VPWR VPWR _4907_/D
+ sky130_fd_sc_hd__o221a_1
X_3209_ _3209_/A VGND VGND VPWR VPWR _3209_/Y sky130_fd_sc_hd__inv_2
X_4189_ _4189_/A VGND VGND VPWR VPWR _4189_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3560_ _5061_/Q _3558_/Y _3488_/B _3559_/X VGND VGND VPWR VPWR _5061_/D sky130_fd_sc_hd__o211a_1
X_2511_ _2519_/A VGND VGND VPWR VPWR _2511_/X sky130_fd_sc_hd__buf_1
X_3491_ input1/X VGND VGND VPWR VPWR _3518_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2442_ _2442_/A VGND VGND VPWR VPWR _2442_/Y sky130_fd_sc_hd__inv_2
X_4112_ _4111_/A _4252_/A _4093_/Y _4094_/X _4111_/X VGND VGND VPWR VPWR _4250_/A
+ sky130_fd_sc_hd__o311a_2
X_5092_ _3386_/X _5092_/D VGND VGND VPWR VPWR _5092_/Q sky130_fd_sc_hd__dfxtp_1
X_4043_ _4886_/Q _4043_/B VGND VGND VPWR VPWR _4043_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4945_ _5018_/CLK _4945_/D VGND VGND VPWR VPWR _4945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4876_ _5028_/CLK _4876_/D VGND VGND VPWR VPWR _4876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3827_ _3827_/A VGND VGND VPWR VPWR _3827_/Y sky130_fd_sc_hd__inv_2
X_3758_ _3758_/A VGND VGND VPWR VPWR _3759_/B sky130_fd_sc_hd__inv_2
X_2709_ _2774_/A VGND VGND VPWR VPWR _2709_/X sky130_fd_sc_hd__buf_1
X_3689_ _3692_/A _3689_/B VGND VGND VPWR VPWR _4997_/D sky130_fd_sc_hd__nor2_1
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2991_ _2991_/A VGND VGND VPWR VPWR _2991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4730_ _4791_/Q _5104_/Q _4729_/Y VGND VGND VPWR VPWR _4731_/A sky130_fd_sc_hd__a21oi_2
X_4661_ _4661_/A VGND VGND VPWR VPWR _4664_/A sky130_fd_sc_hd__inv_2
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3612_ _3612_/A VGND VGND VPWR VPWR _3622_/A sky130_fd_sc_hd__buf_1
X_4592_ _4592_/A _4596_/A VGND VGND VPWR VPWR _4592_/X sky130_fd_sc_hd__or2_1
XFILLER_6_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3543_ _3485_/A _3514_/X _3520_/X _3542_/X VGND VGND VPWR VPWR _3544_/C sky130_fd_sc_hd__a211o_1
X_3474_ _5048_/Q _5049_/Q _5050_/Q VGND VGND VPWR VPWR _3574_/A sky130_fd_sc_hd__and3_1
X_2425_ _2428_/A VGND VGND VPWR VPWR _2425_/X sky130_fd_sc_hd__buf_1
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5075_ _3437_/X _5075_/D VGND VGND VPWR VPWR _5075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4026_ _3673_/B _5004_/Q _3673_/B _5004_/Q VGND VGND VPWR VPWR _4162_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4928_ _5047_/CLK _4928_/D VGND VGND VPWR VPWR _4928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4859_ _5047_/CLK _4859_/D VGND VGND VPWR VPWR _4859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3190_ _3350_/A _2949_/Y _3189_/X VGND VGND VPWR VPWR _3191_/A sky130_fd_sc_hd__o21ai_1
XFILLER_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2974_ _3201_/A _3199_/A VGND VGND VPWR VPWR _2985_/A sky130_fd_sc_hd__nand2_1
X_4713_ _4713_/A VGND VGND VPWR VPWR _4714_/B sky130_fd_sc_hd__inv_2
X_4644_ _4644_/A _4644_/B VGND VGND VPWR VPWR _4828_/D sky130_fd_sc_hd__nor2_1
X_4575_ _4575_/A VGND VGND VPWR VPWR _4575_/X sky130_fd_sc_hd__buf_2
X_3526_ _2899_/X _3518_/A _5048_/Q _3512_/A VGND VGND VPWR VPWR _3531_/A sky130_fd_sc_hd__o22a_1
X_3457_ _5068_/Q _3456_/Y _3435_/X _3457_/C1 VGND VGND VPWR VPWR _5068_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3388_ _5092_/Q _3387_/Y _3375_/X _3388_/C1 VGND VGND VPWR VPWR _5092_/D sky130_fd_sc_hd__o211a_1
X_2408_ _4649_/X _2406_/Y _2407_/Y _2406_/A _4575_/X VGND VGND VPWR VPWR _4824_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5127_ _3204_/X _5127_/D VGND VGND VPWR VPWR _5127_/Q sky130_fd_sc_hd__dfxtp_1
X_5058_ _5063_/CLK _5058_/D VGND VGND VPWR VPWR _5058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4009_ _4899_/Q _5010_/Q _4899_/Q _5010_/Q VGND VGND VPWR VPWR _4010_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2690_ _2690_/A _2690_/B _2690_/C _2690_/D VGND VGND VPWR VPWR _2690_/X sky130_fd_sc_hd__or4_1
XANTENNA_3 _4578_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4360_ _4802_/Q VGND VGND VPWR VPWR _4434_/A sky130_fd_sc_hd__inv_2
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3311_ _3083_/Y _3310_/Y _3083_/A _3310_/A _3267_/X VGND VGND VPWR VPWR _5104_/D
+ sky130_fd_sc_hd__o221a_1
X_4291_ _4291_/A VGND VGND VPWR VPWR _4613_/B sky130_fd_sc_hd__buf_1
X_3242_ _3250_/A _3242_/B VGND VGND VPWR VPWR _3242_/X sky130_fd_sc_hd__or2_1
X_3173_ _3173_/A VGND VGND VPWR VPWR _3173_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer26 _3333_/B VGND VGND VPWR VPWR _3441_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer15 _3349_/B VGND VGND VPWR VPWR _3390_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer37 _3348_/B VGND VGND VPWR VPWR _3392_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer48 _3350_/B VGND VGND VPWR VPWR _3387_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_22_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2957_ _3189_/A _2957_/B VGND VGND VPWR VPWR _2965_/A sky130_fd_sc_hd__or2_1
X_2888_ _2850_/A _3518_/B _3502_/B VGND VGND VPWR VPWR _2889_/A sky130_fd_sc_hd__a21bo_1
X_4627_ _4639_/A VGND VGND VPWR VPWR _4632_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4558_ _4632_/B _4838_/Q _4557_/X VGND VGND VPWR VPWR _4559_/A sky130_fd_sc_hd__o21ai_1
X_4489_ _4517_/A _4320_/X _4460_/X VGND VGND VPWR VPWR _4490_/A sky130_fd_sc_hd__o21ai_2
X_3509_ _3506_/Y _3507_/Y _3508_/X VGND VGND VPWR VPWR _3509_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3860_ _3860_/A _3948_/B VGND VGND VPWR VPWR _3861_/B sky130_fd_sc_hd__or2_1
X_2811_ _2811_/A _2821_/B VGND VGND VPWR VPWR _2811_/X sky130_fd_sc_hd__or2_1
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3791_ _3616_/B _5030_/Q _3618_/B _5029_/Q VGND VGND VPWR VPWR _3791_/X sky130_fd_sc_hd__a211o_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2742_ _2742_/A _2742_/B _2742_/C _2742_/D VGND VGND VPWR VPWR _2745_/B sky130_fd_sc_hd__or4_4
XFILLER_12_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4412_ _4420_/A _4828_/Q _4420_/A _4828_/Q VGND VGND VPWR VPWR _4596_/A sky130_fd_sc_hd__a2bb2o_1
X_2673_ _2703_/A _2624_/B _2590_/D VGND VGND VPWR VPWR _2674_/D sky130_fd_sc_hd__o21a_1
X_4343_ _4805_/Q VGND VGND VPWR VPWR _4343_/X sky130_fd_sc_hd__clkbuf_2
X_4274_ _4863_/Q _4103_/Y _3742_/B _4974_/Q VGND VGND VPWR VPWR _4275_/B sky130_fd_sc_hd__o22a_1
X_3225_ _3225_/A VGND VGND VPWR VPWR _3241_/A sky130_fd_sc_hd__buf_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3156_ _3151_/A _3150_/Y _3151_/Y _3150_/A _3660_/A VGND VGND VPWR VPWR _5137_/D
+ sky130_fd_sc_hd__o221a_1
X_3087_ _3324_/D _3086_/X _5066_/Q _5103_/Q VGND VGND VPWR VPWR _3088_/A sky130_fd_sc_hd__o22a_1
XFILLER_27_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3989_ _3989_/A _3989_/B VGND VGND VPWR VPWR _3989_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer6 _3324_/B VGND VGND VPWR VPWR _3465_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3010_ _3237_/A _3235_/A VGND VGND VPWR VPWR _3125_/A sky130_fd_sc_hd__nand2_1
X_4961_ _5018_/CLK _4961_/D VGND VGND VPWR VPWR _4961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4892_ _5047_/CLK _4892_/D VGND VGND VPWR VPWR _4892_/Q sky130_fd_sc_hd__dfxtp_1
X_3912_ _3923_/A _3775_/B _3870_/Y VGND VGND VPWR VPWR _3913_/B sky130_fd_sc_hd__o21ai_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3843_ _3654_/B _5013_/Q _3833_/Y _3652_/B _5014_/Q VGND VGND VPWR VPWR _3843_/X
+ sky130_fd_sc_hd__o32a_1
X_3774_ _3774_/A _3923_/B VGND VGND VPWR VPWR _3775_/B sky130_fd_sc_hd__or2_1
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2725_ _2680_/A _2705_/X _2693_/X VGND VGND VPWR VPWR _2730_/A sky130_fd_sc_hd__o21a_1
X_2656_ _2656_/A _2656_/B _2656_/C _2656_/D VGND VGND VPWR VPWR _2665_/B sky130_fd_sc_hd__or4_4
X_2587_ _3498_/A _3502_/B _3501_/Y _2587_/D VGND VGND VPWR VPWR _2588_/A sky130_fd_sc_hd__or4_4
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4326_ _4326_/A VGND VGND VPWR VPWR _4620_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4257_ _4257_/A VGND VGND VPWR VPWR _4257_/Y sky130_fd_sc_hd__inv_2
X_4188_ _3687_/B _4998_/Q _4193_/B VGND VGND VPWR VPWR _4189_/A sky130_fd_sc_hd__o21ai_1
X_3208_ _3346_/A _2981_/Y _3207_/X VGND VGND VPWR VPWR _3209_/A sky130_fd_sc_hd__o21ai_1
XFILLER_27_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3139_ _3352_/A _2960_/X _2962_/Y _3353_/A _3138_/Y VGND VGND VPWR VPWR _3139_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_23_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2510_ _4700_/B _2505_/B _2486_/X _2505_/Y VGND VGND VPWR VPWR _4802_/D sky130_fd_sc_hd__o211a_1
X_3490_ input7/X VGND VGND VPWR VPWR _3490_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2441_ _4613_/B _2949_/Y _2440_/X VGND VGND VPWR VPWR _2442_/A sky130_fd_sc_hd__o21ai_1
X_4111_ _4111_/A _4252_/A _4111_/C _4253_/A VGND VGND VPWR VPWR _4111_/X sky130_fd_sc_hd__or4_4
X_5091_ _3389_/X _5091_/D VGND VGND VPWR VPWR _5091_/Q sky130_fd_sc_hd__dfxtp_1
X_4042_ _4997_/Q VGND VGND VPWR VPWR _4043_/B sky130_fd_sc_hd__inv_2
XFILLER_64_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4944_ _5018_/CLK _4944_/D VGND VGND VPWR VPWR _4944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4875_ _5028_/CLK _4875_/D VGND VGND VPWR VPWR _4875_/Q sky130_fd_sc_hd__dfxtp_1
X_3826_ _3824_/A _5016_/Q _3824_/Y _3825_/Y VGND VGND VPWR VPWR _3827_/A sky130_fd_sc_hd__o2bb2a_1
X_3757_ _3593_/B _5040_/Q _4929_/Q _3756_/Y VGND VGND VPWR VPWR _3758_/A sky130_fd_sc_hd__o22a_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2708_ _4941_/Q _2651_/X _2707_/X VGND VGND VPWR VPWR _2715_/B sky130_fd_sc_hd__o21a_1
X_3688_ _4886_/Q VGND VGND VPWR VPWR _3689_/B sky130_fd_sc_hd__inv_2
X_2639_ _4942_/Q _2638_/X _2590_/A VGND VGND VPWR VPWR _2639_/Y sky130_fd_sc_hd__o21ai_1
X_4309_ _4458_/A _4852_/Q _4458_/A _4852_/Q VGND VGND VPWR VPWR _4505_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2990_ _5123_/Q VGND VGND VPWR VPWR _2991_/A sky130_fd_sc_hd__inv_2
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4660_ _4816_/Q _5129_/Q _4291_/A _2949_/Y VGND VGND VPWR VPWR _4661_/A sky130_fd_sc_hd__o22a_1
X_3611_ _3611_/A _3611_/B VGND VGND VPWR VPWR _5032_/D sky130_fd_sc_hd__nor2_1
X_4591_ _4587_/A _4587_/B _4562_/X _4588_/A VGND VGND VPWR VPWR _4867_/D sky130_fd_sc_hd__o211a_1
X_3542_ _3542_/A _3542_/B _3542_/C _3542_/D VGND VGND VPWR VPWR _3542_/X sky130_fd_sc_hd__or4_4
X_3473_ _5058_/Q VGND VGND VPWR VPWR _3484_/A sky130_fd_sc_hd__inv_2
XFILLER_69_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2424_ _4657_/Y _2422_/Y _4657_/A _2422_/A _2423_/X VGND VGND VPWR VPWR _4821_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5074_ _3439_/X _5074_/D VGND VGND VPWR VPWR _5074_/Q sky130_fd_sc_hd__dfxtp_1
X_4025_ _4175_/A _4025_/B VGND VGND VPWR VPWR _4032_/A sky130_fd_sc_hd__or2_1
XFILLER_71_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4927_ _5047_/CLK _4927_/D VGND VGND VPWR VPWR _4927_/Q sky130_fd_sc_hd__dfxtp_1
X_4858_ _5047_/CLK _4858_/D VGND VGND VPWR VPWR _4858_/Q sky130_fd_sc_hd__dfxtp_1
X_3809_ _3809_/A _3809_/B VGND VGND VPWR VPWR _3809_/X sky130_fd_sc_hd__or2_1
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4789_ _2560_/X _4789_/D VGND VGND VPWR VPWR _4789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2973_ _3348_/A _2972_/X _5090_/Q _5127_/Q VGND VGND VPWR VPWR _3199_/A sky130_fd_sc_hd__o22a_1
X_4712_ _4384_/A _3054_/Y _4796_/Q _5109_/Q VGND VGND VPWR VPWR _4713_/A sky130_fd_sc_hd__o22a_1
X_4643_ _4644_/A _4643_/B VGND VGND VPWR VPWR _4829_/D sky130_fd_sc_hd__nor2_1
X_4574_ _4574_/A VGND VGND VPWR VPWR _4574_/Y sky130_fd_sc_hd__inv_2
X_3525_ _3525_/A _3525_/B VGND VGND VPWR VPWR _3525_/Y sky130_fd_sc_hd__nor2_1
X_3456_ _3456_/A VGND VGND VPWR VPWR _3456_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3387_ _3387_/A VGND VGND VPWR VPWR _3387_/Y sky130_fd_sc_hd__clkinvlp_2
X_2407_ _4649_/X VGND VGND VPWR VPWR _2407_/Y sky130_fd_sc_hd__inv_2
X_5126_ _3206_/X _5126_/D VGND VGND VPWR VPWR _5126_/Q sky130_fd_sc_hd__dfxtp_1
X_5057_ _5063_/CLK _5057_/D VGND VGND VPWR VPWR _5057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4008_ _4601_/A _4008_/B VGND VGND VPWR VPWR _4937_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 _4621_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3310_ _3310_/A VGND VGND VPWR VPWR _3310_/Y sky130_fd_sc_hd__inv_2
X_4290_ _4816_/Q VGND VGND VPWR VPWR _4291_/A sky130_fd_sc_hd__inv_2
X_3241_ _3241_/A VGND VGND VPWR VPWR _3241_/X sky130_fd_sc_hd__buf_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3172_ _3172_/A VGND VGND VPWR VPWR _3172_/X sky130_fd_sc_hd__buf_1
XFILLER_66_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer27 _3333_/B VGND VGND VPWR VPWR _3438_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer16 _3341_/B VGND VGND VPWR VPWR _3418_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer38 _3347_/B VGND VGND VPWR VPWR _3398_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer49 _3352_/B VGND VGND VPWR VPWR _3380_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_47_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2956_ _2956_/A VGND VGND VPWR VPWR _2957_/B sky130_fd_sc_hd__inv_2
X_2887_ _5063_/Q _2859_/A _2880_/Y _2922_/C _2886_/X VGND VGND VPWR VPWR _2887_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4626_ _4626_/A _4626_/B VGND VGND VPWR VPWR _4843_/D sky130_fd_sc_hd__nor2_1
X_4557_ _4561_/A _4557_/B VGND VGND VPWR VPWR _4557_/X sky130_fd_sc_hd__or2_1
X_4488_ _4488_/A VGND VGND VPWR VPWR _4492_/A sky130_fd_sc_hd__inv_2
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3508_ _3508_/A _3508_/B VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__or2_1
X_3439_ _3442_/A VGND VGND VPWR VPWR _3439_/X sky130_fd_sc_hd__buf_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5109_ _3285_/X _5109_/D VGND VGND VPWR VPWR _5109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput30 _4777_/Q VGND VGND VPWR VPWR DATA[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2810_ _2810_/A _2810_/B _2810_/C _2810_/D VGND VGND VPWR VPWR _2810_/X sky130_fd_sc_hd__or4_4
X_3790_ _4917_/Q _3787_/Y _3789_/X VGND VGND VPWR VPWR _3790_/Y sky130_fd_sc_hd__o21ai_1
X_2741_ _2768_/A _2712_/X _2713_/X VGND VGND VPWR VPWR _2742_/D sky130_fd_sc_hd__o21a_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4411_ _4790_/Q VGND VGND VPWR VPWR _4420_/A sky130_fd_sc_hd__inv_2
X_2672_ _4950_/Q VGND VGND VPWR VPWR _2703_/A sky130_fd_sc_hd__clkbuf_2
X_4342_ _4342_/A _4534_/A VGND VGND VPWR VPWR _4446_/A sky130_fd_sc_hd__or2_1
X_4273_ _4863_/Q _4103_/Y _4105_/X _3996_/X _4106_/Y VGND VGND VPWR VPWR _4901_/D
+ sky130_fd_sc_hd__o311a_1
X_3224_ _3218_/A _3218_/B _3223_/X _3218_/Y VGND VGND VPWR VPWR _5123_/D sky130_fd_sc_hd__o211a_1
.ends

