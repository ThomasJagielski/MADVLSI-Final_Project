magic
tech sky130A
timestamp 1620315906
<< metal3 >>
rect -115 85 415 515
rect -115 -15 515 85
<< mimcap >>
rect -100 295 400 500
rect -100 205 105 295
rect 195 205 400 295
rect -100 0 400 205
<< mimcapcontact >>
rect 105 205 195 295
<< metal4 >>
rect 100 295 515 300
rect 100 205 105 295
rect 195 205 515 295
rect 100 200 515 205
<< end >>
