magic
tech sky130A
magscale 1 2
timestamp 1620268543
<< pwell >>
rect -4000 1643 -3204 1796
rect -4000 1153 -3847 1643
rect -3357 1153 -3204 1643
rect -4000 1000 -3204 1153
rect -3000 1643 -2204 1796
rect -3000 1153 -2847 1643
rect -2357 1153 -2204 1643
rect -3000 1000 -2204 1153
rect -2000 1643 -1204 1796
rect -2000 1153 -1847 1643
rect -1357 1153 -1204 1643
rect -2000 1000 -1204 1153
rect -1000 1643 -204 1796
rect -1000 1153 -847 1643
rect -357 1153 -204 1643
rect -1000 1000 -204 1153
rect 0 1643 796 1796
rect 0 1153 153 1643
rect 643 1153 796 1643
rect 0 1000 796 1153
rect 1000 1643 1796 1796
rect 1000 1153 1153 1643
rect 1643 1153 1796 1643
rect 1000 1000 1796 1153
rect 2000 1643 2796 1796
rect 2000 1153 2153 1643
rect 2643 1153 2796 1643
rect 2000 1000 2796 1153
rect 3000 1643 3796 1796
rect 3000 1153 3153 1643
rect 3643 1153 3796 1643
rect 3000 1000 3796 1153
rect -4000 643 -3204 796
rect -4000 153 -3847 643
rect -3357 153 -3204 643
rect -4000 0 -3204 153
rect -3000 643 -2204 796
rect -3000 153 -2847 643
rect -2357 153 -2204 643
rect -3000 0 -2204 153
rect -2000 643 -1204 796
rect -2000 153 -1847 643
rect -1357 153 -1204 643
rect -2000 0 -1204 153
rect -1000 643 -204 796
rect -1000 153 -847 643
rect -357 153 -204 643
rect -1000 0 -204 153
rect 1000 643 1796 796
rect 1000 153 1153 643
rect 1643 153 1796 643
rect 1000 0 1796 153
rect 2000 643 2796 796
rect 2000 153 2153 643
rect 2643 153 2796 643
rect 2000 0 2796 153
rect 3000 643 3796 796
rect 3000 153 3153 643
rect 3643 153 3796 643
rect 3000 0 3796 153
rect -4000 -357 -3204 -204
rect -4000 -847 -3847 -357
rect -3357 -847 -3204 -357
rect -4000 -1000 -3204 -847
rect -3000 -357 -2204 -204
rect -3000 -847 -2847 -357
rect -2357 -847 -2204 -357
rect -3000 -1000 -2204 -847
rect -2000 -357 -1204 -204
rect -2000 -847 -1847 -357
rect -1357 -847 -1204 -357
rect -2000 -1000 -1204 -847
rect -1000 -357 -204 -204
rect -1000 -847 -847 -357
rect -357 -847 -204 -357
rect -1000 -1000 -204 -847
rect 0 -357 796 -204
rect 0 -847 153 -357
rect 643 -847 796 -357
rect 0 -1000 796 -847
rect 1000 -357 1796 -204
rect 1000 -847 1153 -357
rect 1643 -847 1796 -357
rect 1000 -1000 1796 -847
rect 2000 -357 2796 -204
rect 2000 -847 2153 -357
rect 2643 -847 2796 -357
rect 2000 -1000 2796 -847
rect 3000 -357 3796 -204
rect 3000 -847 3153 -357
rect 3643 -847 3796 -357
rect 3000 -1000 3796 -847
rect -1000 -1357 -204 -1204
rect -1000 -1847 -847 -1357
rect -357 -1847 -204 -1357
rect -1000 -2000 -204 -1847
rect 0 -1357 796 -1204
rect 0 -1847 153 -1357
rect 643 -1847 796 -1357
rect 0 -2000 796 -1847
rect 1000 -1357 1796 -1204
rect 1000 -1847 1153 -1357
rect 1643 -1847 1796 -1357
rect 1000 -2000 1796 -1847
rect 2000 -1357 2796 -1204
rect 2000 -1847 2153 -1357
rect 2643 -1847 2796 -1357
rect 2000 -2000 2796 -1847
rect 3000 -1357 3796 -1204
rect 3000 -1847 3153 -1357
rect 3643 -1847 3796 -1357
rect 3000 -2000 3796 -1847
rect -1000 -2357 -204 -2204
rect -1000 -2847 -847 -2357
rect -357 -2847 -204 -2357
rect -1000 -3000 -204 -2847
rect 0 -2357 796 -2204
rect 0 -2847 153 -2357
rect 643 -2847 796 -2357
rect 0 -3000 796 -2847
rect 1000 -2357 1796 -2204
rect 1000 -2847 1153 -2357
rect 1643 -2847 1796 -2357
rect 1000 -3000 1796 -2847
rect 2000 -2357 2796 -2204
rect 2000 -2847 2153 -2357
rect 2643 -2847 2796 -2357
rect 2000 -3000 2796 -2847
rect 3000 -2357 3796 -2204
rect 3000 -2847 3153 -2357
rect 3643 -2847 3796 -2357
rect 3000 -3000 3796 -2847
<< nbase >>
rect -3847 1153 -3357 1643
rect -2847 1153 -2357 1643
rect -1847 1153 -1357 1643
rect -847 1153 -357 1643
rect 153 1153 643 1643
rect 1153 1153 1643 1643
rect 2153 1153 2643 1643
rect 3153 1153 3643 1643
rect -3847 153 -3357 643
rect -2847 153 -2357 643
rect -1847 153 -1357 643
rect -847 153 -357 643
rect 1153 153 1643 643
rect 2153 153 2643 643
rect 3153 153 3643 643
rect -3847 -847 -3357 -357
rect -2847 -847 -2357 -357
rect -1847 -847 -1357 -357
rect -847 -847 -357 -357
rect 153 -847 643 -357
rect 1153 -847 1643 -357
rect 2153 -847 2643 -357
rect 3153 -847 3643 -357
rect -847 -1847 -357 -1357
rect 153 -1847 643 -1357
rect 1153 -1847 1643 -1357
rect 2153 -1847 2643 -1357
rect 3153 -1847 3643 -1357
rect -847 -2847 -357 -2357
rect 153 -2847 643 -2357
rect 1153 -2847 1643 -2357
rect 2153 -2847 2643 -2357
rect 3153 -2847 3643 -2357
<< pdiff >>
rect -3670 1449 -3534 1466
rect -3670 1347 -3653 1449
rect -3551 1347 -3534 1449
rect -3670 1330 -3534 1347
rect -2670 1449 -2534 1466
rect -2670 1347 -2653 1449
rect -2551 1347 -2534 1449
rect -2670 1330 -2534 1347
rect -1670 1449 -1534 1466
rect -1670 1347 -1653 1449
rect -1551 1347 -1534 1449
rect -1670 1330 -1534 1347
rect -670 1449 -534 1466
rect -670 1347 -653 1449
rect -551 1347 -534 1449
rect -670 1330 -534 1347
rect 330 1449 466 1466
rect 330 1347 347 1449
rect 449 1347 466 1449
rect 330 1330 466 1347
rect 1330 1449 1466 1466
rect 1330 1347 1347 1449
rect 1449 1347 1466 1449
rect 1330 1330 1466 1347
rect 2330 1449 2466 1466
rect 2330 1347 2347 1449
rect 2449 1347 2466 1449
rect 2330 1330 2466 1347
rect 3330 1449 3466 1466
rect 3330 1347 3347 1449
rect 3449 1347 3466 1449
rect 3330 1330 3466 1347
rect -3670 449 -3534 466
rect -3670 347 -3653 449
rect -3551 347 -3534 449
rect -3670 330 -3534 347
rect -2670 449 -2534 466
rect -2670 347 -2653 449
rect -2551 347 -2534 449
rect -2670 330 -2534 347
rect -1670 449 -1534 466
rect -1670 347 -1653 449
rect -1551 347 -1534 449
rect -1670 330 -1534 347
rect -670 449 -534 466
rect -670 347 -653 449
rect -551 347 -534 449
rect -670 330 -534 347
rect 1330 449 1466 466
rect 1330 347 1347 449
rect 1449 347 1466 449
rect 1330 330 1466 347
rect 2330 449 2466 466
rect 2330 347 2347 449
rect 2449 347 2466 449
rect 2330 330 2466 347
rect 3330 449 3466 466
rect 3330 347 3347 449
rect 3449 347 3466 449
rect 3330 330 3466 347
rect -3670 -551 -3534 -534
rect -3670 -653 -3653 -551
rect -3551 -653 -3534 -551
rect -3670 -670 -3534 -653
rect -2670 -551 -2534 -534
rect -2670 -653 -2653 -551
rect -2551 -653 -2534 -551
rect -2670 -670 -2534 -653
rect -1670 -551 -1534 -534
rect -1670 -653 -1653 -551
rect -1551 -653 -1534 -551
rect -1670 -670 -1534 -653
rect -670 -551 -534 -534
rect -670 -653 -653 -551
rect -551 -653 -534 -551
rect -670 -670 -534 -653
rect 330 -551 466 -534
rect 330 -653 347 -551
rect 449 -653 466 -551
rect 330 -670 466 -653
rect 1330 -551 1466 -534
rect 1330 -653 1347 -551
rect 1449 -653 1466 -551
rect 1330 -670 1466 -653
rect 2330 -551 2466 -534
rect 2330 -653 2347 -551
rect 2449 -653 2466 -551
rect 2330 -670 2466 -653
rect 3330 -551 3466 -534
rect 3330 -653 3347 -551
rect 3449 -653 3466 -551
rect 3330 -670 3466 -653
rect -670 -1551 -534 -1534
rect -670 -1653 -653 -1551
rect -551 -1653 -534 -1551
rect -670 -1670 -534 -1653
rect 330 -1551 466 -1534
rect 330 -1653 347 -1551
rect 449 -1653 466 -1551
rect 330 -1670 466 -1653
rect 1330 -1551 1466 -1534
rect 1330 -1653 1347 -1551
rect 1449 -1653 1466 -1551
rect 1330 -1670 1466 -1653
rect 2330 -1551 2466 -1534
rect 2330 -1653 2347 -1551
rect 2449 -1653 2466 -1551
rect 2330 -1670 2466 -1653
rect 3330 -1551 3466 -1534
rect 3330 -1653 3347 -1551
rect 3449 -1653 3466 -1551
rect 3330 -1670 3466 -1653
rect -670 -2551 -534 -2534
rect -670 -2653 -653 -2551
rect -551 -2653 -534 -2551
rect -670 -2670 -534 -2653
rect 330 -2551 466 -2534
rect 330 -2653 347 -2551
rect 449 -2653 466 -2551
rect 330 -2670 466 -2653
rect 1330 -2551 1466 -2534
rect 1330 -2653 1347 -2551
rect 1449 -2653 1466 -2551
rect 1330 -2670 1466 -2653
rect 2330 -2551 2466 -2534
rect 2330 -2653 2347 -2551
rect 2449 -2653 2466 -2551
rect 2330 -2670 2466 -2653
rect 3330 -2551 3466 -2534
rect 3330 -2653 3347 -2551
rect 3449 -2653 3466 -2551
rect 3330 -2670 3466 -2653
<< pdiffc >>
rect -3653 1347 -3551 1449
rect -2653 1347 -2551 1449
rect -1653 1347 -1551 1449
rect -653 1347 -551 1449
rect 347 1347 449 1449
rect 1347 1347 1449 1449
rect 2347 1347 2449 1449
rect 3347 1347 3449 1449
rect -3653 347 -3551 449
rect -2653 347 -2551 449
rect -1653 347 -1551 449
rect -653 347 -551 449
rect 1347 347 1449 449
rect 2347 347 2449 449
rect 3347 347 3449 449
rect -3653 -653 -3551 -551
rect -2653 -653 -2551 -551
rect -1653 -653 -1551 -551
rect -653 -653 -551 -551
rect 347 -653 449 -551
rect 1347 -653 1449 -551
rect 2347 -653 2449 -551
rect 3347 -653 3449 -551
rect -653 -1653 -551 -1551
rect 347 -1653 449 -1551
rect 1347 -1653 1449 -1551
rect 2347 -1653 2449 -1551
rect 3347 -1653 3449 -1551
rect -653 -2653 -551 -2551
rect 347 -2653 449 -2551
rect 1347 -2653 1449 -2551
rect 2347 -2653 2449 -2551
rect 3347 -2653 3449 -2551
<< psubdiff >>
rect -3974 1736 -3230 1770
rect -3974 1702 -3940 1736
rect -3906 1702 -3872 1736
rect -3838 1702 -3804 1736
rect -3770 1702 -3736 1736
rect -3702 1702 -3502 1736
rect -3468 1702 -3434 1736
rect -3400 1702 -3366 1736
rect -3332 1702 -3298 1736
rect -3264 1702 -3230 1736
rect -3974 1669 -3230 1702
rect -3974 1668 -3873 1669
rect -3974 1634 -3940 1668
rect -3906 1634 -3873 1668
rect -3974 1600 -3873 1634
rect -3331 1668 -3230 1669
rect -3331 1634 -3298 1668
rect -3264 1634 -3230 1668
rect -3974 1566 -3940 1600
rect -3906 1566 -3873 1600
rect -3974 1532 -3873 1566
rect -3974 1498 -3940 1532
rect -3906 1498 -3873 1532
rect -3974 1298 -3873 1498
rect -3974 1264 -3940 1298
rect -3906 1264 -3873 1298
rect -3974 1230 -3873 1264
rect -3974 1196 -3940 1230
rect -3906 1196 -3873 1230
rect -3974 1162 -3873 1196
rect -3331 1600 -3230 1634
rect -3331 1566 -3298 1600
rect -3264 1566 -3230 1600
rect -3331 1532 -3230 1566
rect -3331 1498 -3298 1532
rect -3264 1498 -3230 1532
rect -3331 1298 -3230 1498
rect -3331 1264 -3298 1298
rect -3264 1264 -3230 1298
rect -3331 1230 -3230 1264
rect -3331 1196 -3298 1230
rect -3264 1196 -3230 1230
rect -3974 1128 -3940 1162
rect -3906 1128 -3873 1162
rect -3974 1127 -3873 1128
rect -3331 1162 -3230 1196
rect -3331 1128 -3298 1162
rect -3264 1128 -3230 1162
rect -3331 1127 -3230 1128
rect -3974 1094 -3230 1127
rect -3974 1060 -3940 1094
rect -3906 1060 -3872 1094
rect -3838 1060 -3804 1094
rect -3770 1060 -3736 1094
rect -3702 1060 -3502 1094
rect -3468 1060 -3434 1094
rect -3400 1060 -3366 1094
rect -3332 1060 -3298 1094
rect -3264 1060 -3230 1094
rect -3974 1026 -3230 1060
rect -2974 1736 -2230 1770
rect -2974 1702 -2940 1736
rect -2906 1702 -2872 1736
rect -2838 1702 -2804 1736
rect -2770 1702 -2736 1736
rect -2702 1702 -2502 1736
rect -2468 1702 -2434 1736
rect -2400 1702 -2366 1736
rect -2332 1702 -2298 1736
rect -2264 1702 -2230 1736
rect -2974 1669 -2230 1702
rect -2974 1668 -2873 1669
rect -2974 1634 -2940 1668
rect -2906 1634 -2873 1668
rect -2974 1600 -2873 1634
rect -2331 1668 -2230 1669
rect -2331 1634 -2298 1668
rect -2264 1634 -2230 1668
rect -2974 1566 -2940 1600
rect -2906 1566 -2873 1600
rect -2974 1532 -2873 1566
rect -2974 1498 -2940 1532
rect -2906 1498 -2873 1532
rect -2974 1298 -2873 1498
rect -2974 1264 -2940 1298
rect -2906 1264 -2873 1298
rect -2974 1230 -2873 1264
rect -2974 1196 -2940 1230
rect -2906 1196 -2873 1230
rect -2974 1162 -2873 1196
rect -2331 1600 -2230 1634
rect -2331 1566 -2298 1600
rect -2264 1566 -2230 1600
rect -2331 1532 -2230 1566
rect -2331 1498 -2298 1532
rect -2264 1498 -2230 1532
rect -2331 1298 -2230 1498
rect -2331 1264 -2298 1298
rect -2264 1264 -2230 1298
rect -2331 1230 -2230 1264
rect -2331 1196 -2298 1230
rect -2264 1196 -2230 1230
rect -2974 1128 -2940 1162
rect -2906 1128 -2873 1162
rect -2974 1127 -2873 1128
rect -2331 1162 -2230 1196
rect -2331 1128 -2298 1162
rect -2264 1128 -2230 1162
rect -2331 1127 -2230 1128
rect -2974 1094 -2230 1127
rect -2974 1060 -2940 1094
rect -2906 1060 -2872 1094
rect -2838 1060 -2804 1094
rect -2770 1060 -2736 1094
rect -2702 1060 -2502 1094
rect -2468 1060 -2434 1094
rect -2400 1060 -2366 1094
rect -2332 1060 -2298 1094
rect -2264 1060 -2230 1094
rect -2974 1026 -2230 1060
rect -1974 1736 -1230 1770
rect -1974 1702 -1940 1736
rect -1906 1702 -1872 1736
rect -1838 1702 -1804 1736
rect -1770 1702 -1736 1736
rect -1702 1702 -1502 1736
rect -1468 1702 -1434 1736
rect -1400 1702 -1366 1736
rect -1332 1702 -1298 1736
rect -1264 1702 -1230 1736
rect -1974 1669 -1230 1702
rect -1974 1668 -1873 1669
rect -1974 1634 -1940 1668
rect -1906 1634 -1873 1668
rect -1974 1600 -1873 1634
rect -1331 1668 -1230 1669
rect -1331 1634 -1298 1668
rect -1264 1634 -1230 1668
rect -1974 1566 -1940 1600
rect -1906 1566 -1873 1600
rect -1974 1532 -1873 1566
rect -1974 1498 -1940 1532
rect -1906 1498 -1873 1532
rect -1974 1298 -1873 1498
rect -1974 1264 -1940 1298
rect -1906 1264 -1873 1298
rect -1974 1230 -1873 1264
rect -1974 1196 -1940 1230
rect -1906 1196 -1873 1230
rect -1974 1162 -1873 1196
rect -1331 1600 -1230 1634
rect -1331 1566 -1298 1600
rect -1264 1566 -1230 1600
rect -1331 1532 -1230 1566
rect -1331 1498 -1298 1532
rect -1264 1498 -1230 1532
rect -1331 1298 -1230 1498
rect -1331 1264 -1298 1298
rect -1264 1264 -1230 1298
rect -1331 1230 -1230 1264
rect -1331 1196 -1298 1230
rect -1264 1196 -1230 1230
rect -1974 1128 -1940 1162
rect -1906 1128 -1873 1162
rect -1974 1127 -1873 1128
rect -1331 1162 -1230 1196
rect -1331 1128 -1298 1162
rect -1264 1128 -1230 1162
rect -1331 1127 -1230 1128
rect -1974 1094 -1230 1127
rect -1974 1060 -1940 1094
rect -1906 1060 -1872 1094
rect -1838 1060 -1804 1094
rect -1770 1060 -1736 1094
rect -1702 1060 -1502 1094
rect -1468 1060 -1434 1094
rect -1400 1060 -1366 1094
rect -1332 1060 -1298 1094
rect -1264 1060 -1230 1094
rect -1974 1026 -1230 1060
rect -974 1736 -230 1770
rect -974 1702 -940 1736
rect -906 1702 -872 1736
rect -838 1702 -804 1736
rect -770 1702 -736 1736
rect -702 1702 -502 1736
rect -468 1702 -434 1736
rect -400 1702 -366 1736
rect -332 1702 -298 1736
rect -264 1702 -230 1736
rect -974 1669 -230 1702
rect -974 1668 -873 1669
rect -974 1634 -940 1668
rect -906 1634 -873 1668
rect -974 1600 -873 1634
rect -331 1668 -230 1669
rect -331 1634 -298 1668
rect -264 1634 -230 1668
rect -974 1566 -940 1600
rect -906 1566 -873 1600
rect -974 1532 -873 1566
rect -974 1498 -940 1532
rect -906 1498 -873 1532
rect -974 1298 -873 1498
rect -974 1264 -940 1298
rect -906 1264 -873 1298
rect -974 1230 -873 1264
rect -974 1196 -940 1230
rect -906 1196 -873 1230
rect -974 1162 -873 1196
rect -331 1600 -230 1634
rect -331 1566 -298 1600
rect -264 1566 -230 1600
rect -331 1532 -230 1566
rect -331 1498 -298 1532
rect -264 1498 -230 1532
rect -331 1298 -230 1498
rect -331 1264 -298 1298
rect -264 1264 -230 1298
rect -331 1230 -230 1264
rect -331 1196 -298 1230
rect -264 1196 -230 1230
rect -974 1128 -940 1162
rect -906 1128 -873 1162
rect -974 1127 -873 1128
rect -331 1162 -230 1196
rect -331 1128 -298 1162
rect -264 1128 -230 1162
rect -331 1127 -230 1128
rect -974 1094 -230 1127
rect -974 1060 -940 1094
rect -906 1060 -872 1094
rect -838 1060 -804 1094
rect -770 1060 -736 1094
rect -702 1060 -502 1094
rect -468 1060 -434 1094
rect -400 1060 -366 1094
rect -332 1060 -298 1094
rect -264 1060 -230 1094
rect -974 1026 -230 1060
rect 26 1736 770 1770
rect 26 1702 60 1736
rect 94 1702 128 1736
rect 162 1702 196 1736
rect 230 1702 264 1736
rect 298 1702 498 1736
rect 532 1702 566 1736
rect 600 1702 634 1736
rect 668 1702 702 1736
rect 736 1702 770 1736
rect 26 1669 770 1702
rect 26 1668 127 1669
rect 26 1634 60 1668
rect 94 1634 127 1668
rect 26 1600 127 1634
rect 669 1668 770 1669
rect 669 1634 702 1668
rect 736 1634 770 1668
rect 26 1566 60 1600
rect 94 1566 127 1600
rect 26 1532 127 1566
rect 26 1498 60 1532
rect 94 1498 127 1532
rect 26 1298 127 1498
rect 26 1264 60 1298
rect 94 1264 127 1298
rect 26 1230 127 1264
rect 26 1196 60 1230
rect 94 1196 127 1230
rect 26 1162 127 1196
rect 669 1600 770 1634
rect 669 1566 702 1600
rect 736 1566 770 1600
rect 669 1532 770 1566
rect 669 1498 702 1532
rect 736 1498 770 1532
rect 669 1298 770 1498
rect 669 1264 702 1298
rect 736 1264 770 1298
rect 669 1230 770 1264
rect 669 1196 702 1230
rect 736 1196 770 1230
rect 26 1128 60 1162
rect 94 1128 127 1162
rect 26 1127 127 1128
rect 669 1162 770 1196
rect 669 1128 702 1162
rect 736 1128 770 1162
rect 669 1127 770 1128
rect 26 1094 770 1127
rect 26 1060 60 1094
rect 94 1060 128 1094
rect 162 1060 196 1094
rect 230 1060 264 1094
rect 298 1060 498 1094
rect 532 1060 566 1094
rect 600 1060 634 1094
rect 668 1060 702 1094
rect 736 1060 770 1094
rect 26 1026 770 1060
rect 1026 1736 1770 1770
rect 1026 1702 1060 1736
rect 1094 1702 1128 1736
rect 1162 1702 1196 1736
rect 1230 1702 1264 1736
rect 1298 1702 1498 1736
rect 1532 1702 1566 1736
rect 1600 1702 1634 1736
rect 1668 1702 1702 1736
rect 1736 1702 1770 1736
rect 1026 1669 1770 1702
rect 1026 1668 1127 1669
rect 1026 1634 1060 1668
rect 1094 1634 1127 1668
rect 1026 1600 1127 1634
rect 1669 1668 1770 1669
rect 1669 1634 1702 1668
rect 1736 1634 1770 1668
rect 1026 1566 1060 1600
rect 1094 1566 1127 1600
rect 1026 1532 1127 1566
rect 1026 1498 1060 1532
rect 1094 1498 1127 1532
rect 1026 1298 1127 1498
rect 1026 1264 1060 1298
rect 1094 1264 1127 1298
rect 1026 1230 1127 1264
rect 1026 1196 1060 1230
rect 1094 1196 1127 1230
rect 1026 1162 1127 1196
rect 1669 1600 1770 1634
rect 1669 1566 1702 1600
rect 1736 1566 1770 1600
rect 1669 1532 1770 1566
rect 1669 1498 1702 1532
rect 1736 1498 1770 1532
rect 1669 1298 1770 1498
rect 1669 1264 1702 1298
rect 1736 1264 1770 1298
rect 1669 1230 1770 1264
rect 1669 1196 1702 1230
rect 1736 1196 1770 1230
rect 1026 1128 1060 1162
rect 1094 1128 1127 1162
rect 1026 1127 1127 1128
rect 1669 1162 1770 1196
rect 1669 1128 1702 1162
rect 1736 1128 1770 1162
rect 1669 1127 1770 1128
rect 1026 1094 1770 1127
rect 1026 1060 1060 1094
rect 1094 1060 1128 1094
rect 1162 1060 1196 1094
rect 1230 1060 1264 1094
rect 1298 1060 1498 1094
rect 1532 1060 1566 1094
rect 1600 1060 1634 1094
rect 1668 1060 1702 1094
rect 1736 1060 1770 1094
rect 1026 1026 1770 1060
rect 2026 1736 2770 1770
rect 2026 1702 2060 1736
rect 2094 1702 2128 1736
rect 2162 1702 2196 1736
rect 2230 1702 2264 1736
rect 2298 1702 2498 1736
rect 2532 1702 2566 1736
rect 2600 1702 2634 1736
rect 2668 1702 2702 1736
rect 2736 1702 2770 1736
rect 2026 1669 2770 1702
rect 2026 1668 2127 1669
rect 2026 1634 2060 1668
rect 2094 1634 2127 1668
rect 2026 1600 2127 1634
rect 2669 1668 2770 1669
rect 2669 1634 2702 1668
rect 2736 1634 2770 1668
rect 2026 1566 2060 1600
rect 2094 1566 2127 1600
rect 2026 1532 2127 1566
rect 2026 1498 2060 1532
rect 2094 1498 2127 1532
rect 2026 1298 2127 1498
rect 2026 1264 2060 1298
rect 2094 1264 2127 1298
rect 2026 1230 2127 1264
rect 2026 1196 2060 1230
rect 2094 1196 2127 1230
rect 2026 1162 2127 1196
rect 2669 1600 2770 1634
rect 2669 1566 2702 1600
rect 2736 1566 2770 1600
rect 2669 1532 2770 1566
rect 2669 1498 2702 1532
rect 2736 1498 2770 1532
rect 2669 1298 2770 1498
rect 2669 1264 2702 1298
rect 2736 1264 2770 1298
rect 2669 1230 2770 1264
rect 2669 1196 2702 1230
rect 2736 1196 2770 1230
rect 2026 1128 2060 1162
rect 2094 1128 2127 1162
rect 2026 1127 2127 1128
rect 2669 1162 2770 1196
rect 2669 1128 2702 1162
rect 2736 1128 2770 1162
rect 2669 1127 2770 1128
rect 2026 1094 2770 1127
rect 2026 1060 2060 1094
rect 2094 1060 2128 1094
rect 2162 1060 2196 1094
rect 2230 1060 2264 1094
rect 2298 1060 2498 1094
rect 2532 1060 2566 1094
rect 2600 1060 2634 1094
rect 2668 1060 2702 1094
rect 2736 1060 2770 1094
rect 2026 1026 2770 1060
rect 3026 1736 3770 1770
rect 3026 1702 3060 1736
rect 3094 1702 3128 1736
rect 3162 1702 3196 1736
rect 3230 1702 3264 1736
rect 3298 1702 3498 1736
rect 3532 1702 3566 1736
rect 3600 1702 3634 1736
rect 3668 1702 3702 1736
rect 3736 1702 3770 1736
rect 3026 1669 3770 1702
rect 3026 1668 3127 1669
rect 3026 1634 3060 1668
rect 3094 1634 3127 1668
rect 3026 1600 3127 1634
rect 3669 1668 3770 1669
rect 3669 1634 3702 1668
rect 3736 1634 3770 1668
rect 3026 1566 3060 1600
rect 3094 1566 3127 1600
rect 3026 1532 3127 1566
rect 3026 1498 3060 1532
rect 3094 1498 3127 1532
rect 3026 1298 3127 1498
rect 3026 1264 3060 1298
rect 3094 1264 3127 1298
rect 3026 1230 3127 1264
rect 3026 1196 3060 1230
rect 3094 1196 3127 1230
rect 3026 1162 3127 1196
rect 3669 1600 3770 1634
rect 3669 1566 3702 1600
rect 3736 1566 3770 1600
rect 3669 1532 3770 1566
rect 3669 1498 3702 1532
rect 3736 1498 3770 1532
rect 3669 1298 3770 1498
rect 3669 1264 3702 1298
rect 3736 1264 3770 1298
rect 3669 1230 3770 1264
rect 3669 1196 3702 1230
rect 3736 1196 3770 1230
rect 3026 1128 3060 1162
rect 3094 1128 3127 1162
rect 3026 1127 3127 1128
rect 3669 1162 3770 1196
rect 3669 1128 3702 1162
rect 3736 1128 3770 1162
rect 3669 1127 3770 1128
rect 3026 1094 3770 1127
rect 3026 1060 3060 1094
rect 3094 1060 3128 1094
rect 3162 1060 3196 1094
rect 3230 1060 3264 1094
rect 3298 1060 3498 1094
rect 3532 1060 3566 1094
rect 3600 1060 3634 1094
rect 3668 1060 3702 1094
rect 3736 1060 3770 1094
rect 3026 1026 3770 1060
rect -3974 736 -3230 770
rect -3974 702 -3940 736
rect -3906 702 -3872 736
rect -3838 702 -3804 736
rect -3770 702 -3736 736
rect -3702 702 -3502 736
rect -3468 702 -3434 736
rect -3400 702 -3366 736
rect -3332 702 -3298 736
rect -3264 702 -3230 736
rect -3974 669 -3230 702
rect -3974 668 -3873 669
rect -3974 634 -3940 668
rect -3906 634 -3873 668
rect -3974 600 -3873 634
rect -3331 668 -3230 669
rect -3331 634 -3298 668
rect -3264 634 -3230 668
rect -3974 566 -3940 600
rect -3906 566 -3873 600
rect -3974 532 -3873 566
rect -3974 498 -3940 532
rect -3906 498 -3873 532
rect -3974 298 -3873 498
rect -3974 264 -3940 298
rect -3906 264 -3873 298
rect -3974 230 -3873 264
rect -3974 196 -3940 230
rect -3906 196 -3873 230
rect -3974 162 -3873 196
rect -3331 600 -3230 634
rect -3331 566 -3298 600
rect -3264 566 -3230 600
rect -3331 532 -3230 566
rect -3331 498 -3298 532
rect -3264 498 -3230 532
rect -3331 298 -3230 498
rect -3331 264 -3298 298
rect -3264 264 -3230 298
rect -3331 230 -3230 264
rect -3331 196 -3298 230
rect -3264 196 -3230 230
rect -3974 128 -3940 162
rect -3906 128 -3873 162
rect -3974 127 -3873 128
rect -3331 162 -3230 196
rect -3331 128 -3298 162
rect -3264 128 -3230 162
rect -3331 127 -3230 128
rect -3974 94 -3230 127
rect -3974 60 -3940 94
rect -3906 60 -3872 94
rect -3838 60 -3804 94
rect -3770 60 -3736 94
rect -3702 60 -3502 94
rect -3468 60 -3434 94
rect -3400 60 -3366 94
rect -3332 60 -3298 94
rect -3264 60 -3230 94
rect -3974 26 -3230 60
rect -2974 736 -2230 770
rect -2974 702 -2940 736
rect -2906 702 -2872 736
rect -2838 702 -2804 736
rect -2770 702 -2736 736
rect -2702 702 -2502 736
rect -2468 702 -2434 736
rect -2400 702 -2366 736
rect -2332 702 -2298 736
rect -2264 702 -2230 736
rect -2974 669 -2230 702
rect -2974 668 -2873 669
rect -2974 634 -2940 668
rect -2906 634 -2873 668
rect -2974 600 -2873 634
rect -2331 668 -2230 669
rect -2331 634 -2298 668
rect -2264 634 -2230 668
rect -2974 566 -2940 600
rect -2906 566 -2873 600
rect -2974 532 -2873 566
rect -2974 498 -2940 532
rect -2906 498 -2873 532
rect -2974 298 -2873 498
rect -2974 264 -2940 298
rect -2906 264 -2873 298
rect -2974 230 -2873 264
rect -2974 196 -2940 230
rect -2906 196 -2873 230
rect -2974 162 -2873 196
rect -2331 600 -2230 634
rect -2331 566 -2298 600
rect -2264 566 -2230 600
rect -2331 532 -2230 566
rect -2331 498 -2298 532
rect -2264 498 -2230 532
rect -2331 298 -2230 498
rect -2331 264 -2298 298
rect -2264 264 -2230 298
rect -2331 230 -2230 264
rect -2331 196 -2298 230
rect -2264 196 -2230 230
rect -2974 128 -2940 162
rect -2906 128 -2873 162
rect -2974 127 -2873 128
rect -2331 162 -2230 196
rect -2331 128 -2298 162
rect -2264 128 -2230 162
rect -2331 127 -2230 128
rect -2974 94 -2230 127
rect -2974 60 -2940 94
rect -2906 60 -2872 94
rect -2838 60 -2804 94
rect -2770 60 -2736 94
rect -2702 60 -2502 94
rect -2468 60 -2434 94
rect -2400 60 -2366 94
rect -2332 60 -2298 94
rect -2264 60 -2230 94
rect -2974 26 -2230 60
rect -1974 736 -1230 770
rect -1974 702 -1940 736
rect -1906 702 -1872 736
rect -1838 702 -1804 736
rect -1770 702 -1736 736
rect -1702 702 -1502 736
rect -1468 702 -1434 736
rect -1400 702 -1366 736
rect -1332 702 -1298 736
rect -1264 702 -1230 736
rect -1974 669 -1230 702
rect -1974 668 -1873 669
rect -1974 634 -1940 668
rect -1906 634 -1873 668
rect -1974 600 -1873 634
rect -1331 668 -1230 669
rect -1331 634 -1298 668
rect -1264 634 -1230 668
rect -1974 566 -1940 600
rect -1906 566 -1873 600
rect -1974 532 -1873 566
rect -1974 498 -1940 532
rect -1906 498 -1873 532
rect -1974 298 -1873 498
rect -1974 264 -1940 298
rect -1906 264 -1873 298
rect -1974 230 -1873 264
rect -1974 196 -1940 230
rect -1906 196 -1873 230
rect -1974 162 -1873 196
rect -1331 600 -1230 634
rect -1331 566 -1298 600
rect -1264 566 -1230 600
rect -1331 532 -1230 566
rect -1331 498 -1298 532
rect -1264 498 -1230 532
rect -1331 298 -1230 498
rect -1331 264 -1298 298
rect -1264 264 -1230 298
rect -1331 230 -1230 264
rect -1331 196 -1298 230
rect -1264 196 -1230 230
rect -1974 128 -1940 162
rect -1906 128 -1873 162
rect -1974 127 -1873 128
rect -1331 162 -1230 196
rect -1331 128 -1298 162
rect -1264 128 -1230 162
rect -1331 127 -1230 128
rect -1974 94 -1230 127
rect -1974 60 -1940 94
rect -1906 60 -1872 94
rect -1838 60 -1804 94
rect -1770 60 -1736 94
rect -1702 60 -1502 94
rect -1468 60 -1434 94
rect -1400 60 -1366 94
rect -1332 60 -1298 94
rect -1264 60 -1230 94
rect -1974 26 -1230 60
rect -974 736 -230 770
rect -974 702 -940 736
rect -906 702 -872 736
rect -838 702 -804 736
rect -770 702 -736 736
rect -702 702 -502 736
rect -468 702 -434 736
rect -400 702 -366 736
rect -332 702 -298 736
rect -264 702 -230 736
rect -974 669 -230 702
rect -974 668 -873 669
rect -974 634 -940 668
rect -906 634 -873 668
rect -974 600 -873 634
rect -331 668 -230 669
rect -331 634 -298 668
rect -264 634 -230 668
rect -974 566 -940 600
rect -906 566 -873 600
rect -974 532 -873 566
rect -974 498 -940 532
rect -906 498 -873 532
rect -974 298 -873 498
rect -974 264 -940 298
rect -906 264 -873 298
rect -974 230 -873 264
rect -974 196 -940 230
rect -906 196 -873 230
rect -974 162 -873 196
rect -331 600 -230 634
rect -331 566 -298 600
rect -264 566 -230 600
rect -331 532 -230 566
rect -331 498 -298 532
rect -264 498 -230 532
rect -331 298 -230 498
rect -331 264 -298 298
rect -264 264 -230 298
rect -331 230 -230 264
rect -331 196 -298 230
rect -264 196 -230 230
rect -974 128 -940 162
rect -906 128 -873 162
rect -974 127 -873 128
rect -331 162 -230 196
rect -331 128 -298 162
rect -264 128 -230 162
rect -331 127 -230 128
rect -974 94 -230 127
rect -974 60 -940 94
rect -906 60 -872 94
rect -838 60 -804 94
rect -770 60 -736 94
rect -702 60 -502 94
rect -468 60 -434 94
rect -400 60 -366 94
rect -332 60 -298 94
rect -264 60 -230 94
rect -974 26 -230 60
rect 1026 736 1770 770
rect 1026 702 1060 736
rect 1094 702 1128 736
rect 1162 702 1196 736
rect 1230 702 1264 736
rect 1298 702 1498 736
rect 1532 702 1566 736
rect 1600 702 1634 736
rect 1668 702 1702 736
rect 1736 702 1770 736
rect 1026 669 1770 702
rect 1026 668 1127 669
rect 1026 634 1060 668
rect 1094 634 1127 668
rect 1026 600 1127 634
rect 1669 668 1770 669
rect 1669 634 1702 668
rect 1736 634 1770 668
rect 1026 566 1060 600
rect 1094 566 1127 600
rect 1026 532 1127 566
rect 1026 498 1060 532
rect 1094 498 1127 532
rect 1026 298 1127 498
rect 1026 264 1060 298
rect 1094 264 1127 298
rect 1026 230 1127 264
rect 1026 196 1060 230
rect 1094 196 1127 230
rect 1026 162 1127 196
rect 1669 600 1770 634
rect 1669 566 1702 600
rect 1736 566 1770 600
rect 1669 532 1770 566
rect 1669 498 1702 532
rect 1736 498 1770 532
rect 1669 298 1770 498
rect 1669 264 1702 298
rect 1736 264 1770 298
rect 1669 230 1770 264
rect 1669 196 1702 230
rect 1736 196 1770 230
rect 1026 128 1060 162
rect 1094 128 1127 162
rect 1026 127 1127 128
rect 1669 162 1770 196
rect 1669 128 1702 162
rect 1736 128 1770 162
rect 1669 127 1770 128
rect 1026 94 1770 127
rect 1026 60 1060 94
rect 1094 60 1128 94
rect 1162 60 1196 94
rect 1230 60 1264 94
rect 1298 60 1498 94
rect 1532 60 1566 94
rect 1600 60 1634 94
rect 1668 60 1702 94
rect 1736 60 1770 94
rect 1026 26 1770 60
rect 2026 736 2770 770
rect 2026 702 2060 736
rect 2094 702 2128 736
rect 2162 702 2196 736
rect 2230 702 2264 736
rect 2298 702 2498 736
rect 2532 702 2566 736
rect 2600 702 2634 736
rect 2668 702 2702 736
rect 2736 702 2770 736
rect 2026 669 2770 702
rect 2026 668 2127 669
rect 2026 634 2060 668
rect 2094 634 2127 668
rect 2026 600 2127 634
rect 2669 668 2770 669
rect 2669 634 2702 668
rect 2736 634 2770 668
rect 2026 566 2060 600
rect 2094 566 2127 600
rect 2026 532 2127 566
rect 2026 498 2060 532
rect 2094 498 2127 532
rect 2026 298 2127 498
rect 2026 264 2060 298
rect 2094 264 2127 298
rect 2026 230 2127 264
rect 2026 196 2060 230
rect 2094 196 2127 230
rect 2026 162 2127 196
rect 2669 600 2770 634
rect 2669 566 2702 600
rect 2736 566 2770 600
rect 2669 532 2770 566
rect 2669 498 2702 532
rect 2736 498 2770 532
rect 2669 298 2770 498
rect 2669 264 2702 298
rect 2736 264 2770 298
rect 2669 230 2770 264
rect 2669 196 2702 230
rect 2736 196 2770 230
rect 2026 128 2060 162
rect 2094 128 2127 162
rect 2026 127 2127 128
rect 2669 162 2770 196
rect 2669 128 2702 162
rect 2736 128 2770 162
rect 2669 127 2770 128
rect 2026 94 2770 127
rect 2026 60 2060 94
rect 2094 60 2128 94
rect 2162 60 2196 94
rect 2230 60 2264 94
rect 2298 60 2498 94
rect 2532 60 2566 94
rect 2600 60 2634 94
rect 2668 60 2702 94
rect 2736 60 2770 94
rect 2026 26 2770 60
rect 3026 736 3770 770
rect 3026 702 3060 736
rect 3094 702 3128 736
rect 3162 702 3196 736
rect 3230 702 3264 736
rect 3298 702 3498 736
rect 3532 702 3566 736
rect 3600 702 3634 736
rect 3668 702 3702 736
rect 3736 702 3770 736
rect 3026 669 3770 702
rect 3026 668 3127 669
rect 3026 634 3060 668
rect 3094 634 3127 668
rect 3026 600 3127 634
rect 3669 668 3770 669
rect 3669 634 3702 668
rect 3736 634 3770 668
rect 3026 566 3060 600
rect 3094 566 3127 600
rect 3026 532 3127 566
rect 3026 498 3060 532
rect 3094 498 3127 532
rect 3026 298 3127 498
rect 3026 264 3060 298
rect 3094 264 3127 298
rect 3026 230 3127 264
rect 3026 196 3060 230
rect 3094 196 3127 230
rect 3026 162 3127 196
rect 3669 600 3770 634
rect 3669 566 3702 600
rect 3736 566 3770 600
rect 3669 532 3770 566
rect 3669 498 3702 532
rect 3736 498 3770 532
rect 3669 298 3770 498
rect 3669 264 3702 298
rect 3736 264 3770 298
rect 3669 230 3770 264
rect 3669 196 3702 230
rect 3736 196 3770 230
rect 3026 128 3060 162
rect 3094 128 3127 162
rect 3026 127 3127 128
rect 3669 162 3770 196
rect 3669 128 3702 162
rect 3736 128 3770 162
rect 3669 127 3770 128
rect 3026 94 3770 127
rect 3026 60 3060 94
rect 3094 60 3128 94
rect 3162 60 3196 94
rect 3230 60 3264 94
rect 3298 60 3498 94
rect 3532 60 3566 94
rect 3600 60 3634 94
rect 3668 60 3702 94
rect 3736 60 3770 94
rect 3026 26 3770 60
rect -3974 -264 -3230 -230
rect -3974 -298 -3940 -264
rect -3906 -298 -3872 -264
rect -3838 -298 -3804 -264
rect -3770 -298 -3736 -264
rect -3702 -298 -3502 -264
rect -3468 -298 -3434 -264
rect -3400 -298 -3366 -264
rect -3332 -298 -3298 -264
rect -3264 -298 -3230 -264
rect -3974 -331 -3230 -298
rect -3974 -332 -3873 -331
rect -3974 -366 -3940 -332
rect -3906 -366 -3873 -332
rect -3974 -400 -3873 -366
rect -3331 -332 -3230 -331
rect -3331 -366 -3298 -332
rect -3264 -366 -3230 -332
rect -3974 -434 -3940 -400
rect -3906 -434 -3873 -400
rect -3974 -468 -3873 -434
rect -3974 -502 -3940 -468
rect -3906 -502 -3873 -468
rect -3974 -702 -3873 -502
rect -3974 -736 -3940 -702
rect -3906 -736 -3873 -702
rect -3974 -770 -3873 -736
rect -3974 -804 -3940 -770
rect -3906 -804 -3873 -770
rect -3974 -838 -3873 -804
rect -3331 -400 -3230 -366
rect -3331 -434 -3298 -400
rect -3264 -434 -3230 -400
rect -3331 -468 -3230 -434
rect -3331 -502 -3298 -468
rect -3264 -502 -3230 -468
rect -3331 -702 -3230 -502
rect -3331 -736 -3298 -702
rect -3264 -736 -3230 -702
rect -3331 -770 -3230 -736
rect -3331 -804 -3298 -770
rect -3264 -804 -3230 -770
rect -3974 -872 -3940 -838
rect -3906 -872 -3873 -838
rect -3974 -873 -3873 -872
rect -3331 -838 -3230 -804
rect -3331 -872 -3298 -838
rect -3264 -872 -3230 -838
rect -3331 -873 -3230 -872
rect -3974 -906 -3230 -873
rect -3974 -940 -3940 -906
rect -3906 -940 -3872 -906
rect -3838 -940 -3804 -906
rect -3770 -940 -3736 -906
rect -3702 -940 -3502 -906
rect -3468 -940 -3434 -906
rect -3400 -940 -3366 -906
rect -3332 -940 -3298 -906
rect -3264 -940 -3230 -906
rect -3974 -974 -3230 -940
rect -2974 -264 -2230 -230
rect -2974 -298 -2940 -264
rect -2906 -298 -2872 -264
rect -2838 -298 -2804 -264
rect -2770 -298 -2736 -264
rect -2702 -298 -2502 -264
rect -2468 -298 -2434 -264
rect -2400 -298 -2366 -264
rect -2332 -298 -2298 -264
rect -2264 -298 -2230 -264
rect -2974 -331 -2230 -298
rect -2974 -332 -2873 -331
rect -2974 -366 -2940 -332
rect -2906 -366 -2873 -332
rect -2974 -400 -2873 -366
rect -2331 -332 -2230 -331
rect -2331 -366 -2298 -332
rect -2264 -366 -2230 -332
rect -2974 -434 -2940 -400
rect -2906 -434 -2873 -400
rect -2974 -468 -2873 -434
rect -2974 -502 -2940 -468
rect -2906 -502 -2873 -468
rect -2974 -702 -2873 -502
rect -2974 -736 -2940 -702
rect -2906 -736 -2873 -702
rect -2974 -770 -2873 -736
rect -2974 -804 -2940 -770
rect -2906 -804 -2873 -770
rect -2974 -838 -2873 -804
rect -2331 -400 -2230 -366
rect -2331 -434 -2298 -400
rect -2264 -434 -2230 -400
rect -2331 -468 -2230 -434
rect -2331 -502 -2298 -468
rect -2264 -502 -2230 -468
rect -2331 -702 -2230 -502
rect -2331 -736 -2298 -702
rect -2264 -736 -2230 -702
rect -2331 -770 -2230 -736
rect -2331 -804 -2298 -770
rect -2264 -804 -2230 -770
rect -2974 -872 -2940 -838
rect -2906 -872 -2873 -838
rect -2974 -873 -2873 -872
rect -2331 -838 -2230 -804
rect -2331 -872 -2298 -838
rect -2264 -872 -2230 -838
rect -2331 -873 -2230 -872
rect -2974 -906 -2230 -873
rect -2974 -940 -2940 -906
rect -2906 -940 -2872 -906
rect -2838 -940 -2804 -906
rect -2770 -940 -2736 -906
rect -2702 -940 -2502 -906
rect -2468 -940 -2434 -906
rect -2400 -940 -2366 -906
rect -2332 -940 -2298 -906
rect -2264 -940 -2230 -906
rect -2974 -974 -2230 -940
rect -1974 -264 -1230 -230
rect -1974 -298 -1940 -264
rect -1906 -298 -1872 -264
rect -1838 -298 -1804 -264
rect -1770 -298 -1736 -264
rect -1702 -298 -1502 -264
rect -1468 -298 -1434 -264
rect -1400 -298 -1366 -264
rect -1332 -298 -1298 -264
rect -1264 -298 -1230 -264
rect -1974 -331 -1230 -298
rect -1974 -332 -1873 -331
rect -1974 -366 -1940 -332
rect -1906 -366 -1873 -332
rect -1974 -400 -1873 -366
rect -1331 -332 -1230 -331
rect -1331 -366 -1298 -332
rect -1264 -366 -1230 -332
rect -1974 -434 -1940 -400
rect -1906 -434 -1873 -400
rect -1974 -468 -1873 -434
rect -1974 -502 -1940 -468
rect -1906 -502 -1873 -468
rect -1974 -702 -1873 -502
rect -1974 -736 -1940 -702
rect -1906 -736 -1873 -702
rect -1974 -770 -1873 -736
rect -1974 -804 -1940 -770
rect -1906 -804 -1873 -770
rect -1974 -838 -1873 -804
rect -1331 -400 -1230 -366
rect -1331 -434 -1298 -400
rect -1264 -434 -1230 -400
rect -1331 -468 -1230 -434
rect -1331 -502 -1298 -468
rect -1264 -502 -1230 -468
rect -1331 -702 -1230 -502
rect -1331 -736 -1298 -702
rect -1264 -736 -1230 -702
rect -1331 -770 -1230 -736
rect -1331 -804 -1298 -770
rect -1264 -804 -1230 -770
rect -1974 -872 -1940 -838
rect -1906 -872 -1873 -838
rect -1974 -873 -1873 -872
rect -1331 -838 -1230 -804
rect -1331 -872 -1298 -838
rect -1264 -872 -1230 -838
rect -1331 -873 -1230 -872
rect -1974 -906 -1230 -873
rect -1974 -940 -1940 -906
rect -1906 -940 -1872 -906
rect -1838 -940 -1804 -906
rect -1770 -940 -1736 -906
rect -1702 -940 -1502 -906
rect -1468 -940 -1434 -906
rect -1400 -940 -1366 -906
rect -1332 -940 -1298 -906
rect -1264 -940 -1230 -906
rect -1974 -974 -1230 -940
rect -974 -264 -230 -230
rect -974 -298 -940 -264
rect -906 -298 -872 -264
rect -838 -298 -804 -264
rect -770 -298 -736 -264
rect -702 -298 -502 -264
rect -468 -298 -434 -264
rect -400 -298 -366 -264
rect -332 -298 -298 -264
rect -264 -298 -230 -264
rect -974 -331 -230 -298
rect -974 -332 -873 -331
rect -974 -366 -940 -332
rect -906 -366 -873 -332
rect -974 -400 -873 -366
rect -331 -332 -230 -331
rect -331 -366 -298 -332
rect -264 -366 -230 -332
rect -974 -434 -940 -400
rect -906 -434 -873 -400
rect -974 -468 -873 -434
rect -974 -502 -940 -468
rect -906 -502 -873 -468
rect -974 -702 -873 -502
rect -974 -736 -940 -702
rect -906 -736 -873 -702
rect -974 -770 -873 -736
rect -974 -804 -940 -770
rect -906 -804 -873 -770
rect -974 -838 -873 -804
rect -331 -400 -230 -366
rect -331 -434 -298 -400
rect -264 -434 -230 -400
rect -331 -468 -230 -434
rect -331 -502 -298 -468
rect -264 -502 -230 -468
rect -331 -702 -230 -502
rect -331 -736 -298 -702
rect -264 -736 -230 -702
rect -331 -770 -230 -736
rect -331 -804 -298 -770
rect -264 -804 -230 -770
rect -974 -872 -940 -838
rect -906 -872 -873 -838
rect -974 -873 -873 -872
rect -331 -838 -230 -804
rect -331 -872 -298 -838
rect -264 -872 -230 -838
rect -331 -873 -230 -872
rect -974 -906 -230 -873
rect -974 -940 -940 -906
rect -906 -940 -872 -906
rect -838 -940 -804 -906
rect -770 -940 -736 -906
rect -702 -940 -502 -906
rect -468 -940 -434 -906
rect -400 -940 -366 -906
rect -332 -940 -298 -906
rect -264 -940 -230 -906
rect -974 -974 -230 -940
rect 26 -264 770 -230
rect 26 -298 60 -264
rect 94 -298 128 -264
rect 162 -298 196 -264
rect 230 -298 264 -264
rect 298 -298 498 -264
rect 532 -298 566 -264
rect 600 -298 634 -264
rect 668 -298 702 -264
rect 736 -298 770 -264
rect 26 -331 770 -298
rect 26 -332 127 -331
rect 26 -366 60 -332
rect 94 -366 127 -332
rect 26 -400 127 -366
rect 669 -332 770 -331
rect 669 -366 702 -332
rect 736 -366 770 -332
rect 26 -434 60 -400
rect 94 -434 127 -400
rect 26 -468 127 -434
rect 26 -502 60 -468
rect 94 -502 127 -468
rect 26 -702 127 -502
rect 26 -736 60 -702
rect 94 -736 127 -702
rect 26 -770 127 -736
rect 26 -804 60 -770
rect 94 -804 127 -770
rect 26 -838 127 -804
rect 669 -400 770 -366
rect 669 -434 702 -400
rect 736 -434 770 -400
rect 669 -468 770 -434
rect 669 -502 702 -468
rect 736 -502 770 -468
rect 669 -702 770 -502
rect 669 -736 702 -702
rect 736 -736 770 -702
rect 669 -770 770 -736
rect 669 -804 702 -770
rect 736 -804 770 -770
rect 26 -872 60 -838
rect 94 -872 127 -838
rect 26 -873 127 -872
rect 669 -838 770 -804
rect 669 -872 702 -838
rect 736 -872 770 -838
rect 669 -873 770 -872
rect 26 -906 770 -873
rect 26 -940 60 -906
rect 94 -940 128 -906
rect 162 -940 196 -906
rect 230 -940 264 -906
rect 298 -940 498 -906
rect 532 -940 566 -906
rect 600 -940 634 -906
rect 668 -940 702 -906
rect 736 -940 770 -906
rect 26 -974 770 -940
rect 1026 -264 1770 -230
rect 1026 -298 1060 -264
rect 1094 -298 1128 -264
rect 1162 -298 1196 -264
rect 1230 -298 1264 -264
rect 1298 -298 1498 -264
rect 1532 -298 1566 -264
rect 1600 -298 1634 -264
rect 1668 -298 1702 -264
rect 1736 -298 1770 -264
rect 1026 -331 1770 -298
rect 1026 -332 1127 -331
rect 1026 -366 1060 -332
rect 1094 -366 1127 -332
rect 1026 -400 1127 -366
rect 1669 -332 1770 -331
rect 1669 -366 1702 -332
rect 1736 -366 1770 -332
rect 1026 -434 1060 -400
rect 1094 -434 1127 -400
rect 1026 -468 1127 -434
rect 1026 -502 1060 -468
rect 1094 -502 1127 -468
rect 1026 -702 1127 -502
rect 1026 -736 1060 -702
rect 1094 -736 1127 -702
rect 1026 -770 1127 -736
rect 1026 -804 1060 -770
rect 1094 -804 1127 -770
rect 1026 -838 1127 -804
rect 1669 -400 1770 -366
rect 1669 -434 1702 -400
rect 1736 -434 1770 -400
rect 1669 -468 1770 -434
rect 1669 -502 1702 -468
rect 1736 -502 1770 -468
rect 1669 -702 1770 -502
rect 1669 -736 1702 -702
rect 1736 -736 1770 -702
rect 1669 -770 1770 -736
rect 1669 -804 1702 -770
rect 1736 -804 1770 -770
rect 1026 -872 1060 -838
rect 1094 -872 1127 -838
rect 1026 -873 1127 -872
rect 1669 -838 1770 -804
rect 1669 -872 1702 -838
rect 1736 -872 1770 -838
rect 1669 -873 1770 -872
rect 1026 -906 1770 -873
rect 1026 -940 1060 -906
rect 1094 -940 1128 -906
rect 1162 -940 1196 -906
rect 1230 -940 1264 -906
rect 1298 -940 1498 -906
rect 1532 -940 1566 -906
rect 1600 -940 1634 -906
rect 1668 -940 1702 -906
rect 1736 -940 1770 -906
rect 1026 -974 1770 -940
rect 2026 -264 2770 -230
rect 2026 -298 2060 -264
rect 2094 -298 2128 -264
rect 2162 -298 2196 -264
rect 2230 -298 2264 -264
rect 2298 -298 2498 -264
rect 2532 -298 2566 -264
rect 2600 -298 2634 -264
rect 2668 -298 2702 -264
rect 2736 -298 2770 -264
rect 2026 -331 2770 -298
rect 2026 -332 2127 -331
rect 2026 -366 2060 -332
rect 2094 -366 2127 -332
rect 2026 -400 2127 -366
rect 2669 -332 2770 -331
rect 2669 -366 2702 -332
rect 2736 -366 2770 -332
rect 2026 -434 2060 -400
rect 2094 -434 2127 -400
rect 2026 -468 2127 -434
rect 2026 -502 2060 -468
rect 2094 -502 2127 -468
rect 2026 -702 2127 -502
rect 2026 -736 2060 -702
rect 2094 -736 2127 -702
rect 2026 -770 2127 -736
rect 2026 -804 2060 -770
rect 2094 -804 2127 -770
rect 2026 -838 2127 -804
rect 2669 -400 2770 -366
rect 2669 -434 2702 -400
rect 2736 -434 2770 -400
rect 2669 -468 2770 -434
rect 2669 -502 2702 -468
rect 2736 -502 2770 -468
rect 2669 -702 2770 -502
rect 2669 -736 2702 -702
rect 2736 -736 2770 -702
rect 2669 -770 2770 -736
rect 2669 -804 2702 -770
rect 2736 -804 2770 -770
rect 2026 -872 2060 -838
rect 2094 -872 2127 -838
rect 2026 -873 2127 -872
rect 2669 -838 2770 -804
rect 2669 -872 2702 -838
rect 2736 -872 2770 -838
rect 2669 -873 2770 -872
rect 2026 -906 2770 -873
rect 2026 -940 2060 -906
rect 2094 -940 2128 -906
rect 2162 -940 2196 -906
rect 2230 -940 2264 -906
rect 2298 -940 2498 -906
rect 2532 -940 2566 -906
rect 2600 -940 2634 -906
rect 2668 -940 2702 -906
rect 2736 -940 2770 -906
rect 2026 -974 2770 -940
rect 3026 -264 3770 -230
rect 3026 -298 3060 -264
rect 3094 -298 3128 -264
rect 3162 -298 3196 -264
rect 3230 -298 3264 -264
rect 3298 -298 3498 -264
rect 3532 -298 3566 -264
rect 3600 -298 3634 -264
rect 3668 -298 3702 -264
rect 3736 -298 3770 -264
rect 3026 -331 3770 -298
rect 3026 -332 3127 -331
rect 3026 -366 3060 -332
rect 3094 -366 3127 -332
rect 3026 -400 3127 -366
rect 3669 -332 3770 -331
rect 3669 -366 3702 -332
rect 3736 -366 3770 -332
rect 3026 -434 3060 -400
rect 3094 -434 3127 -400
rect 3026 -468 3127 -434
rect 3026 -502 3060 -468
rect 3094 -502 3127 -468
rect 3026 -702 3127 -502
rect 3026 -736 3060 -702
rect 3094 -736 3127 -702
rect 3026 -770 3127 -736
rect 3026 -804 3060 -770
rect 3094 -804 3127 -770
rect 3026 -838 3127 -804
rect 3669 -400 3770 -366
rect 3669 -434 3702 -400
rect 3736 -434 3770 -400
rect 3669 -468 3770 -434
rect 3669 -502 3702 -468
rect 3736 -502 3770 -468
rect 3669 -702 3770 -502
rect 3669 -736 3702 -702
rect 3736 -736 3770 -702
rect 3669 -770 3770 -736
rect 3669 -804 3702 -770
rect 3736 -804 3770 -770
rect 3026 -872 3060 -838
rect 3094 -872 3127 -838
rect 3026 -873 3127 -872
rect 3669 -838 3770 -804
rect 3669 -872 3702 -838
rect 3736 -872 3770 -838
rect 3669 -873 3770 -872
rect 3026 -906 3770 -873
rect 3026 -940 3060 -906
rect 3094 -940 3128 -906
rect 3162 -940 3196 -906
rect 3230 -940 3264 -906
rect 3298 -940 3498 -906
rect 3532 -940 3566 -906
rect 3600 -940 3634 -906
rect 3668 -940 3702 -906
rect 3736 -940 3770 -906
rect 3026 -974 3770 -940
rect -974 -1264 -230 -1230
rect -974 -1298 -940 -1264
rect -906 -1298 -872 -1264
rect -838 -1298 -804 -1264
rect -770 -1298 -736 -1264
rect -702 -1298 -502 -1264
rect -468 -1298 -434 -1264
rect -400 -1298 -366 -1264
rect -332 -1298 -298 -1264
rect -264 -1298 -230 -1264
rect -974 -1331 -230 -1298
rect -974 -1332 -873 -1331
rect -974 -1366 -940 -1332
rect -906 -1366 -873 -1332
rect -974 -1400 -873 -1366
rect -331 -1332 -230 -1331
rect -331 -1366 -298 -1332
rect -264 -1366 -230 -1332
rect -974 -1434 -940 -1400
rect -906 -1434 -873 -1400
rect -974 -1468 -873 -1434
rect -974 -1502 -940 -1468
rect -906 -1502 -873 -1468
rect -974 -1702 -873 -1502
rect -974 -1736 -940 -1702
rect -906 -1736 -873 -1702
rect -974 -1770 -873 -1736
rect -974 -1804 -940 -1770
rect -906 -1804 -873 -1770
rect -974 -1838 -873 -1804
rect -331 -1400 -230 -1366
rect -331 -1434 -298 -1400
rect -264 -1434 -230 -1400
rect -331 -1468 -230 -1434
rect -331 -1502 -298 -1468
rect -264 -1502 -230 -1468
rect -331 -1702 -230 -1502
rect -331 -1736 -298 -1702
rect -264 -1736 -230 -1702
rect -331 -1770 -230 -1736
rect -331 -1804 -298 -1770
rect -264 -1804 -230 -1770
rect -974 -1872 -940 -1838
rect -906 -1872 -873 -1838
rect -974 -1873 -873 -1872
rect -331 -1838 -230 -1804
rect -331 -1872 -298 -1838
rect -264 -1872 -230 -1838
rect -331 -1873 -230 -1872
rect -974 -1906 -230 -1873
rect -974 -1940 -940 -1906
rect -906 -1940 -872 -1906
rect -838 -1940 -804 -1906
rect -770 -1940 -736 -1906
rect -702 -1940 -502 -1906
rect -468 -1940 -434 -1906
rect -400 -1940 -366 -1906
rect -332 -1940 -298 -1906
rect -264 -1940 -230 -1906
rect -974 -1974 -230 -1940
rect 26 -1264 770 -1230
rect 26 -1298 60 -1264
rect 94 -1298 128 -1264
rect 162 -1298 196 -1264
rect 230 -1298 264 -1264
rect 298 -1298 498 -1264
rect 532 -1298 566 -1264
rect 600 -1298 634 -1264
rect 668 -1298 702 -1264
rect 736 -1298 770 -1264
rect 26 -1331 770 -1298
rect 26 -1332 127 -1331
rect 26 -1366 60 -1332
rect 94 -1366 127 -1332
rect 26 -1400 127 -1366
rect 669 -1332 770 -1331
rect 669 -1366 702 -1332
rect 736 -1366 770 -1332
rect 26 -1434 60 -1400
rect 94 -1434 127 -1400
rect 26 -1468 127 -1434
rect 26 -1502 60 -1468
rect 94 -1502 127 -1468
rect 26 -1702 127 -1502
rect 26 -1736 60 -1702
rect 94 -1736 127 -1702
rect 26 -1770 127 -1736
rect 26 -1804 60 -1770
rect 94 -1804 127 -1770
rect 26 -1838 127 -1804
rect 669 -1400 770 -1366
rect 669 -1434 702 -1400
rect 736 -1434 770 -1400
rect 669 -1468 770 -1434
rect 669 -1502 702 -1468
rect 736 -1502 770 -1468
rect 669 -1702 770 -1502
rect 669 -1736 702 -1702
rect 736 -1736 770 -1702
rect 669 -1770 770 -1736
rect 669 -1804 702 -1770
rect 736 -1804 770 -1770
rect 26 -1872 60 -1838
rect 94 -1872 127 -1838
rect 26 -1873 127 -1872
rect 669 -1838 770 -1804
rect 669 -1872 702 -1838
rect 736 -1872 770 -1838
rect 669 -1873 770 -1872
rect 26 -1906 770 -1873
rect 26 -1940 60 -1906
rect 94 -1940 128 -1906
rect 162 -1940 196 -1906
rect 230 -1940 264 -1906
rect 298 -1940 498 -1906
rect 532 -1940 566 -1906
rect 600 -1940 634 -1906
rect 668 -1940 702 -1906
rect 736 -1940 770 -1906
rect 26 -1974 770 -1940
rect 1026 -1264 1770 -1230
rect 1026 -1298 1060 -1264
rect 1094 -1298 1128 -1264
rect 1162 -1298 1196 -1264
rect 1230 -1298 1264 -1264
rect 1298 -1298 1498 -1264
rect 1532 -1298 1566 -1264
rect 1600 -1298 1634 -1264
rect 1668 -1298 1702 -1264
rect 1736 -1298 1770 -1264
rect 1026 -1331 1770 -1298
rect 1026 -1332 1127 -1331
rect 1026 -1366 1060 -1332
rect 1094 -1366 1127 -1332
rect 1026 -1400 1127 -1366
rect 1669 -1332 1770 -1331
rect 1669 -1366 1702 -1332
rect 1736 -1366 1770 -1332
rect 1026 -1434 1060 -1400
rect 1094 -1434 1127 -1400
rect 1026 -1468 1127 -1434
rect 1026 -1502 1060 -1468
rect 1094 -1502 1127 -1468
rect 1026 -1702 1127 -1502
rect 1026 -1736 1060 -1702
rect 1094 -1736 1127 -1702
rect 1026 -1770 1127 -1736
rect 1026 -1804 1060 -1770
rect 1094 -1804 1127 -1770
rect 1026 -1838 1127 -1804
rect 1669 -1400 1770 -1366
rect 1669 -1434 1702 -1400
rect 1736 -1434 1770 -1400
rect 1669 -1468 1770 -1434
rect 1669 -1502 1702 -1468
rect 1736 -1502 1770 -1468
rect 1669 -1702 1770 -1502
rect 1669 -1736 1702 -1702
rect 1736 -1736 1770 -1702
rect 1669 -1770 1770 -1736
rect 1669 -1804 1702 -1770
rect 1736 -1804 1770 -1770
rect 1026 -1872 1060 -1838
rect 1094 -1872 1127 -1838
rect 1026 -1873 1127 -1872
rect 1669 -1838 1770 -1804
rect 1669 -1872 1702 -1838
rect 1736 -1872 1770 -1838
rect 1669 -1873 1770 -1872
rect 1026 -1906 1770 -1873
rect 1026 -1940 1060 -1906
rect 1094 -1940 1128 -1906
rect 1162 -1940 1196 -1906
rect 1230 -1940 1264 -1906
rect 1298 -1940 1498 -1906
rect 1532 -1940 1566 -1906
rect 1600 -1940 1634 -1906
rect 1668 -1940 1702 -1906
rect 1736 -1940 1770 -1906
rect 1026 -1974 1770 -1940
rect 2026 -1264 2770 -1230
rect 2026 -1298 2060 -1264
rect 2094 -1298 2128 -1264
rect 2162 -1298 2196 -1264
rect 2230 -1298 2264 -1264
rect 2298 -1298 2498 -1264
rect 2532 -1298 2566 -1264
rect 2600 -1298 2634 -1264
rect 2668 -1298 2702 -1264
rect 2736 -1298 2770 -1264
rect 2026 -1331 2770 -1298
rect 2026 -1332 2127 -1331
rect 2026 -1366 2060 -1332
rect 2094 -1366 2127 -1332
rect 2026 -1400 2127 -1366
rect 2669 -1332 2770 -1331
rect 2669 -1366 2702 -1332
rect 2736 -1366 2770 -1332
rect 2026 -1434 2060 -1400
rect 2094 -1434 2127 -1400
rect 2026 -1468 2127 -1434
rect 2026 -1502 2060 -1468
rect 2094 -1502 2127 -1468
rect 2026 -1702 2127 -1502
rect 2026 -1736 2060 -1702
rect 2094 -1736 2127 -1702
rect 2026 -1770 2127 -1736
rect 2026 -1804 2060 -1770
rect 2094 -1804 2127 -1770
rect 2026 -1838 2127 -1804
rect 2669 -1400 2770 -1366
rect 2669 -1434 2702 -1400
rect 2736 -1434 2770 -1400
rect 2669 -1468 2770 -1434
rect 2669 -1502 2702 -1468
rect 2736 -1502 2770 -1468
rect 2669 -1702 2770 -1502
rect 2669 -1736 2702 -1702
rect 2736 -1736 2770 -1702
rect 2669 -1770 2770 -1736
rect 2669 -1804 2702 -1770
rect 2736 -1804 2770 -1770
rect 2026 -1872 2060 -1838
rect 2094 -1872 2127 -1838
rect 2026 -1873 2127 -1872
rect 2669 -1838 2770 -1804
rect 2669 -1872 2702 -1838
rect 2736 -1872 2770 -1838
rect 2669 -1873 2770 -1872
rect 2026 -1906 2770 -1873
rect 2026 -1940 2060 -1906
rect 2094 -1940 2128 -1906
rect 2162 -1940 2196 -1906
rect 2230 -1940 2264 -1906
rect 2298 -1940 2498 -1906
rect 2532 -1940 2566 -1906
rect 2600 -1940 2634 -1906
rect 2668 -1940 2702 -1906
rect 2736 -1940 2770 -1906
rect 2026 -1974 2770 -1940
rect 3026 -1264 3770 -1230
rect 3026 -1298 3060 -1264
rect 3094 -1298 3128 -1264
rect 3162 -1298 3196 -1264
rect 3230 -1298 3264 -1264
rect 3298 -1298 3498 -1264
rect 3532 -1298 3566 -1264
rect 3600 -1298 3634 -1264
rect 3668 -1298 3702 -1264
rect 3736 -1298 3770 -1264
rect 3026 -1331 3770 -1298
rect 3026 -1332 3127 -1331
rect 3026 -1366 3060 -1332
rect 3094 -1366 3127 -1332
rect 3026 -1400 3127 -1366
rect 3669 -1332 3770 -1331
rect 3669 -1366 3702 -1332
rect 3736 -1366 3770 -1332
rect 3026 -1434 3060 -1400
rect 3094 -1434 3127 -1400
rect 3026 -1468 3127 -1434
rect 3026 -1502 3060 -1468
rect 3094 -1502 3127 -1468
rect 3026 -1702 3127 -1502
rect 3026 -1736 3060 -1702
rect 3094 -1736 3127 -1702
rect 3026 -1770 3127 -1736
rect 3026 -1804 3060 -1770
rect 3094 -1804 3127 -1770
rect 3026 -1838 3127 -1804
rect 3669 -1400 3770 -1366
rect 3669 -1434 3702 -1400
rect 3736 -1434 3770 -1400
rect 3669 -1468 3770 -1434
rect 3669 -1502 3702 -1468
rect 3736 -1502 3770 -1468
rect 3669 -1702 3770 -1502
rect 3669 -1736 3702 -1702
rect 3736 -1736 3770 -1702
rect 3669 -1770 3770 -1736
rect 3669 -1804 3702 -1770
rect 3736 -1804 3770 -1770
rect 3026 -1872 3060 -1838
rect 3094 -1872 3127 -1838
rect 3026 -1873 3127 -1872
rect 3669 -1838 3770 -1804
rect 3669 -1872 3702 -1838
rect 3736 -1872 3770 -1838
rect 3669 -1873 3770 -1872
rect 3026 -1906 3770 -1873
rect 3026 -1940 3060 -1906
rect 3094 -1940 3128 -1906
rect 3162 -1940 3196 -1906
rect 3230 -1940 3264 -1906
rect 3298 -1940 3498 -1906
rect 3532 -1940 3566 -1906
rect 3600 -1940 3634 -1906
rect 3668 -1940 3702 -1906
rect 3736 -1940 3770 -1906
rect 3026 -1974 3770 -1940
rect -974 -2264 -230 -2230
rect -974 -2298 -940 -2264
rect -906 -2298 -872 -2264
rect -838 -2298 -804 -2264
rect -770 -2298 -736 -2264
rect -702 -2298 -502 -2264
rect -468 -2298 -434 -2264
rect -400 -2298 -366 -2264
rect -332 -2298 -298 -2264
rect -264 -2298 -230 -2264
rect -974 -2331 -230 -2298
rect -974 -2332 -873 -2331
rect -974 -2366 -940 -2332
rect -906 -2366 -873 -2332
rect -974 -2400 -873 -2366
rect -331 -2332 -230 -2331
rect -331 -2366 -298 -2332
rect -264 -2366 -230 -2332
rect -974 -2434 -940 -2400
rect -906 -2434 -873 -2400
rect -974 -2468 -873 -2434
rect -974 -2502 -940 -2468
rect -906 -2502 -873 -2468
rect -974 -2702 -873 -2502
rect -974 -2736 -940 -2702
rect -906 -2736 -873 -2702
rect -974 -2770 -873 -2736
rect -974 -2804 -940 -2770
rect -906 -2804 -873 -2770
rect -974 -2838 -873 -2804
rect -331 -2400 -230 -2366
rect -331 -2434 -298 -2400
rect -264 -2434 -230 -2400
rect -331 -2468 -230 -2434
rect -331 -2502 -298 -2468
rect -264 -2502 -230 -2468
rect -331 -2702 -230 -2502
rect -331 -2736 -298 -2702
rect -264 -2736 -230 -2702
rect -331 -2770 -230 -2736
rect -331 -2804 -298 -2770
rect -264 -2804 -230 -2770
rect -974 -2872 -940 -2838
rect -906 -2872 -873 -2838
rect -974 -2873 -873 -2872
rect -331 -2838 -230 -2804
rect -331 -2872 -298 -2838
rect -264 -2872 -230 -2838
rect -331 -2873 -230 -2872
rect -974 -2906 -230 -2873
rect -974 -2940 -940 -2906
rect -906 -2940 -872 -2906
rect -838 -2940 -804 -2906
rect -770 -2940 -736 -2906
rect -702 -2940 -502 -2906
rect -468 -2940 -434 -2906
rect -400 -2940 -366 -2906
rect -332 -2940 -298 -2906
rect -264 -2940 -230 -2906
rect -974 -2974 -230 -2940
rect 26 -2264 770 -2230
rect 26 -2298 60 -2264
rect 94 -2298 128 -2264
rect 162 -2298 196 -2264
rect 230 -2298 264 -2264
rect 298 -2298 498 -2264
rect 532 -2298 566 -2264
rect 600 -2298 634 -2264
rect 668 -2298 702 -2264
rect 736 -2298 770 -2264
rect 26 -2331 770 -2298
rect 26 -2332 127 -2331
rect 26 -2366 60 -2332
rect 94 -2366 127 -2332
rect 26 -2400 127 -2366
rect 669 -2332 770 -2331
rect 669 -2366 702 -2332
rect 736 -2366 770 -2332
rect 26 -2434 60 -2400
rect 94 -2434 127 -2400
rect 26 -2468 127 -2434
rect 26 -2502 60 -2468
rect 94 -2502 127 -2468
rect 26 -2702 127 -2502
rect 26 -2736 60 -2702
rect 94 -2736 127 -2702
rect 26 -2770 127 -2736
rect 26 -2804 60 -2770
rect 94 -2804 127 -2770
rect 26 -2838 127 -2804
rect 669 -2400 770 -2366
rect 669 -2434 702 -2400
rect 736 -2434 770 -2400
rect 669 -2468 770 -2434
rect 669 -2502 702 -2468
rect 736 -2502 770 -2468
rect 669 -2702 770 -2502
rect 669 -2736 702 -2702
rect 736 -2736 770 -2702
rect 669 -2770 770 -2736
rect 669 -2804 702 -2770
rect 736 -2804 770 -2770
rect 26 -2872 60 -2838
rect 94 -2872 127 -2838
rect 26 -2873 127 -2872
rect 669 -2838 770 -2804
rect 669 -2872 702 -2838
rect 736 -2872 770 -2838
rect 669 -2873 770 -2872
rect 26 -2906 770 -2873
rect 26 -2940 60 -2906
rect 94 -2940 128 -2906
rect 162 -2940 196 -2906
rect 230 -2940 264 -2906
rect 298 -2940 498 -2906
rect 532 -2940 566 -2906
rect 600 -2940 634 -2906
rect 668 -2940 702 -2906
rect 736 -2940 770 -2906
rect 26 -2974 770 -2940
rect 1026 -2264 1770 -2230
rect 1026 -2298 1060 -2264
rect 1094 -2298 1128 -2264
rect 1162 -2298 1196 -2264
rect 1230 -2298 1264 -2264
rect 1298 -2298 1498 -2264
rect 1532 -2298 1566 -2264
rect 1600 -2298 1634 -2264
rect 1668 -2298 1702 -2264
rect 1736 -2298 1770 -2264
rect 1026 -2331 1770 -2298
rect 1026 -2332 1127 -2331
rect 1026 -2366 1060 -2332
rect 1094 -2366 1127 -2332
rect 1026 -2400 1127 -2366
rect 1669 -2332 1770 -2331
rect 1669 -2366 1702 -2332
rect 1736 -2366 1770 -2332
rect 1026 -2434 1060 -2400
rect 1094 -2434 1127 -2400
rect 1026 -2468 1127 -2434
rect 1026 -2502 1060 -2468
rect 1094 -2502 1127 -2468
rect 1026 -2702 1127 -2502
rect 1026 -2736 1060 -2702
rect 1094 -2736 1127 -2702
rect 1026 -2770 1127 -2736
rect 1026 -2804 1060 -2770
rect 1094 -2804 1127 -2770
rect 1026 -2838 1127 -2804
rect 1669 -2400 1770 -2366
rect 1669 -2434 1702 -2400
rect 1736 -2434 1770 -2400
rect 1669 -2468 1770 -2434
rect 1669 -2502 1702 -2468
rect 1736 -2502 1770 -2468
rect 1669 -2702 1770 -2502
rect 1669 -2736 1702 -2702
rect 1736 -2736 1770 -2702
rect 1669 -2770 1770 -2736
rect 1669 -2804 1702 -2770
rect 1736 -2804 1770 -2770
rect 1026 -2872 1060 -2838
rect 1094 -2872 1127 -2838
rect 1026 -2873 1127 -2872
rect 1669 -2838 1770 -2804
rect 1669 -2872 1702 -2838
rect 1736 -2872 1770 -2838
rect 1669 -2873 1770 -2872
rect 1026 -2906 1770 -2873
rect 1026 -2940 1060 -2906
rect 1094 -2940 1128 -2906
rect 1162 -2940 1196 -2906
rect 1230 -2940 1264 -2906
rect 1298 -2940 1498 -2906
rect 1532 -2940 1566 -2906
rect 1600 -2940 1634 -2906
rect 1668 -2940 1702 -2906
rect 1736 -2940 1770 -2906
rect 1026 -2974 1770 -2940
rect 2026 -2264 2770 -2230
rect 2026 -2298 2060 -2264
rect 2094 -2298 2128 -2264
rect 2162 -2298 2196 -2264
rect 2230 -2298 2264 -2264
rect 2298 -2298 2498 -2264
rect 2532 -2298 2566 -2264
rect 2600 -2298 2634 -2264
rect 2668 -2298 2702 -2264
rect 2736 -2298 2770 -2264
rect 2026 -2331 2770 -2298
rect 2026 -2332 2127 -2331
rect 2026 -2366 2060 -2332
rect 2094 -2366 2127 -2332
rect 2026 -2400 2127 -2366
rect 2669 -2332 2770 -2331
rect 2669 -2366 2702 -2332
rect 2736 -2366 2770 -2332
rect 2026 -2434 2060 -2400
rect 2094 -2434 2127 -2400
rect 2026 -2468 2127 -2434
rect 2026 -2502 2060 -2468
rect 2094 -2502 2127 -2468
rect 2026 -2702 2127 -2502
rect 2026 -2736 2060 -2702
rect 2094 -2736 2127 -2702
rect 2026 -2770 2127 -2736
rect 2026 -2804 2060 -2770
rect 2094 -2804 2127 -2770
rect 2026 -2838 2127 -2804
rect 2669 -2400 2770 -2366
rect 2669 -2434 2702 -2400
rect 2736 -2434 2770 -2400
rect 2669 -2468 2770 -2434
rect 2669 -2502 2702 -2468
rect 2736 -2502 2770 -2468
rect 2669 -2702 2770 -2502
rect 2669 -2736 2702 -2702
rect 2736 -2736 2770 -2702
rect 2669 -2770 2770 -2736
rect 2669 -2804 2702 -2770
rect 2736 -2804 2770 -2770
rect 2026 -2872 2060 -2838
rect 2094 -2872 2127 -2838
rect 2026 -2873 2127 -2872
rect 2669 -2838 2770 -2804
rect 2669 -2872 2702 -2838
rect 2736 -2872 2770 -2838
rect 2669 -2873 2770 -2872
rect 2026 -2906 2770 -2873
rect 2026 -2940 2060 -2906
rect 2094 -2940 2128 -2906
rect 2162 -2940 2196 -2906
rect 2230 -2940 2264 -2906
rect 2298 -2940 2498 -2906
rect 2532 -2940 2566 -2906
rect 2600 -2940 2634 -2906
rect 2668 -2940 2702 -2906
rect 2736 -2940 2770 -2906
rect 2026 -2974 2770 -2940
rect 3026 -2264 3770 -2230
rect 3026 -2298 3060 -2264
rect 3094 -2298 3128 -2264
rect 3162 -2298 3196 -2264
rect 3230 -2298 3264 -2264
rect 3298 -2298 3498 -2264
rect 3532 -2298 3566 -2264
rect 3600 -2298 3634 -2264
rect 3668 -2298 3702 -2264
rect 3736 -2298 3770 -2264
rect 3026 -2331 3770 -2298
rect 3026 -2332 3127 -2331
rect 3026 -2366 3060 -2332
rect 3094 -2366 3127 -2332
rect 3026 -2400 3127 -2366
rect 3669 -2332 3770 -2331
rect 3669 -2366 3702 -2332
rect 3736 -2366 3770 -2332
rect 3026 -2434 3060 -2400
rect 3094 -2434 3127 -2400
rect 3026 -2468 3127 -2434
rect 3026 -2502 3060 -2468
rect 3094 -2502 3127 -2468
rect 3026 -2702 3127 -2502
rect 3026 -2736 3060 -2702
rect 3094 -2736 3127 -2702
rect 3026 -2770 3127 -2736
rect 3026 -2804 3060 -2770
rect 3094 -2804 3127 -2770
rect 3026 -2838 3127 -2804
rect 3669 -2400 3770 -2366
rect 3669 -2434 3702 -2400
rect 3736 -2434 3770 -2400
rect 3669 -2468 3770 -2434
rect 3669 -2502 3702 -2468
rect 3736 -2502 3770 -2468
rect 3669 -2702 3770 -2502
rect 3669 -2736 3702 -2702
rect 3736 -2736 3770 -2702
rect 3669 -2770 3770 -2736
rect 3669 -2804 3702 -2770
rect 3736 -2804 3770 -2770
rect 3026 -2872 3060 -2838
rect 3094 -2872 3127 -2838
rect 3026 -2873 3127 -2872
rect 3669 -2838 3770 -2804
rect 3669 -2872 3702 -2838
rect 3736 -2872 3770 -2838
rect 3669 -2873 3770 -2872
rect 3026 -2906 3770 -2873
rect 3026 -2940 3060 -2906
rect 3094 -2940 3128 -2906
rect 3162 -2940 3196 -2906
rect 3230 -2940 3264 -2906
rect 3298 -2940 3498 -2906
rect 3532 -2940 3566 -2906
rect 3600 -2940 3634 -2906
rect 3668 -2940 3702 -2906
rect 3736 -2940 3770 -2906
rect 3026 -2974 3770 -2940
<< nsubdiff >>
rect -3811 1583 -3393 1607
rect -3811 1549 -3787 1583
rect -3753 1549 -3719 1583
rect -3685 1549 -3519 1583
rect -3485 1549 -3451 1583
rect -3417 1549 -3393 1583
rect -3811 1535 -3393 1549
rect -3811 1515 -3739 1535
rect -3811 1481 -3787 1515
rect -3753 1481 -3739 1515
rect -3811 1315 -3739 1481
rect -3465 1515 -3393 1535
rect -3465 1481 -3451 1515
rect -3417 1481 -3393 1515
rect -3811 1281 -3787 1315
rect -3753 1281 -3739 1315
rect -3811 1261 -3739 1281
rect -3465 1315 -3393 1481
rect -3465 1281 -3451 1315
rect -3417 1281 -3393 1315
rect -3465 1261 -3393 1281
rect -3811 1247 -3393 1261
rect -3811 1213 -3787 1247
rect -3753 1213 -3719 1247
rect -3685 1213 -3519 1247
rect -3485 1213 -3451 1247
rect -3417 1213 -3393 1247
rect -3811 1189 -3393 1213
rect -2811 1583 -2393 1607
rect -2811 1549 -2787 1583
rect -2753 1549 -2719 1583
rect -2685 1549 -2519 1583
rect -2485 1549 -2451 1583
rect -2417 1549 -2393 1583
rect -2811 1535 -2393 1549
rect -2811 1515 -2739 1535
rect -2811 1481 -2787 1515
rect -2753 1481 -2739 1515
rect -2811 1315 -2739 1481
rect -2465 1515 -2393 1535
rect -2465 1481 -2451 1515
rect -2417 1481 -2393 1515
rect -2811 1281 -2787 1315
rect -2753 1281 -2739 1315
rect -2811 1261 -2739 1281
rect -2465 1315 -2393 1481
rect -2465 1281 -2451 1315
rect -2417 1281 -2393 1315
rect -2465 1261 -2393 1281
rect -2811 1247 -2393 1261
rect -2811 1213 -2787 1247
rect -2753 1213 -2719 1247
rect -2685 1213 -2519 1247
rect -2485 1213 -2451 1247
rect -2417 1213 -2393 1247
rect -2811 1189 -2393 1213
rect -1811 1583 -1393 1607
rect -1811 1549 -1787 1583
rect -1753 1549 -1719 1583
rect -1685 1549 -1519 1583
rect -1485 1549 -1451 1583
rect -1417 1549 -1393 1583
rect -1811 1535 -1393 1549
rect -1811 1515 -1739 1535
rect -1811 1481 -1787 1515
rect -1753 1481 -1739 1515
rect -1811 1315 -1739 1481
rect -1465 1515 -1393 1535
rect -1465 1481 -1451 1515
rect -1417 1481 -1393 1515
rect -1811 1281 -1787 1315
rect -1753 1281 -1739 1315
rect -1811 1261 -1739 1281
rect -1465 1315 -1393 1481
rect -1465 1281 -1451 1315
rect -1417 1281 -1393 1315
rect -1465 1261 -1393 1281
rect -1811 1247 -1393 1261
rect -1811 1213 -1787 1247
rect -1753 1213 -1719 1247
rect -1685 1213 -1519 1247
rect -1485 1213 -1451 1247
rect -1417 1213 -1393 1247
rect -1811 1189 -1393 1213
rect -811 1583 -393 1607
rect -811 1549 -787 1583
rect -753 1549 -719 1583
rect -685 1549 -519 1583
rect -485 1549 -451 1583
rect -417 1549 -393 1583
rect -811 1535 -393 1549
rect -811 1515 -739 1535
rect -811 1481 -787 1515
rect -753 1481 -739 1515
rect -811 1315 -739 1481
rect -465 1515 -393 1535
rect -465 1481 -451 1515
rect -417 1481 -393 1515
rect -811 1281 -787 1315
rect -753 1281 -739 1315
rect -811 1261 -739 1281
rect -465 1315 -393 1481
rect -465 1281 -451 1315
rect -417 1281 -393 1315
rect -465 1261 -393 1281
rect -811 1247 -393 1261
rect -811 1213 -787 1247
rect -753 1213 -719 1247
rect -685 1213 -519 1247
rect -485 1213 -451 1247
rect -417 1213 -393 1247
rect -811 1189 -393 1213
rect 189 1583 607 1607
rect 189 1549 213 1583
rect 247 1549 281 1583
rect 315 1549 481 1583
rect 515 1549 549 1583
rect 583 1549 607 1583
rect 189 1535 607 1549
rect 189 1515 261 1535
rect 189 1481 213 1515
rect 247 1481 261 1515
rect 189 1315 261 1481
rect 535 1515 607 1535
rect 535 1481 549 1515
rect 583 1481 607 1515
rect 189 1281 213 1315
rect 247 1281 261 1315
rect 189 1261 261 1281
rect 535 1315 607 1481
rect 535 1281 549 1315
rect 583 1281 607 1315
rect 535 1261 607 1281
rect 189 1247 607 1261
rect 189 1213 213 1247
rect 247 1213 281 1247
rect 315 1213 481 1247
rect 515 1213 549 1247
rect 583 1213 607 1247
rect 189 1189 607 1213
rect 1189 1583 1607 1607
rect 1189 1549 1213 1583
rect 1247 1549 1281 1583
rect 1315 1549 1481 1583
rect 1515 1549 1549 1583
rect 1583 1549 1607 1583
rect 1189 1535 1607 1549
rect 1189 1515 1261 1535
rect 1189 1481 1213 1515
rect 1247 1481 1261 1515
rect 1189 1315 1261 1481
rect 1535 1515 1607 1535
rect 1535 1481 1549 1515
rect 1583 1481 1607 1515
rect 1189 1281 1213 1315
rect 1247 1281 1261 1315
rect 1189 1261 1261 1281
rect 1535 1315 1607 1481
rect 1535 1281 1549 1315
rect 1583 1281 1607 1315
rect 1535 1261 1607 1281
rect 1189 1247 1607 1261
rect 1189 1213 1213 1247
rect 1247 1213 1281 1247
rect 1315 1213 1481 1247
rect 1515 1213 1549 1247
rect 1583 1213 1607 1247
rect 1189 1189 1607 1213
rect 2189 1583 2607 1607
rect 2189 1549 2213 1583
rect 2247 1549 2281 1583
rect 2315 1549 2481 1583
rect 2515 1549 2549 1583
rect 2583 1549 2607 1583
rect 2189 1535 2607 1549
rect 2189 1515 2261 1535
rect 2189 1481 2213 1515
rect 2247 1481 2261 1515
rect 2189 1315 2261 1481
rect 2535 1515 2607 1535
rect 2535 1481 2549 1515
rect 2583 1481 2607 1515
rect 2189 1281 2213 1315
rect 2247 1281 2261 1315
rect 2189 1261 2261 1281
rect 2535 1315 2607 1481
rect 2535 1281 2549 1315
rect 2583 1281 2607 1315
rect 2535 1261 2607 1281
rect 2189 1247 2607 1261
rect 2189 1213 2213 1247
rect 2247 1213 2281 1247
rect 2315 1213 2481 1247
rect 2515 1213 2549 1247
rect 2583 1213 2607 1247
rect 2189 1189 2607 1213
rect 3189 1583 3607 1607
rect 3189 1549 3213 1583
rect 3247 1549 3281 1583
rect 3315 1549 3481 1583
rect 3515 1549 3549 1583
rect 3583 1549 3607 1583
rect 3189 1535 3607 1549
rect 3189 1515 3261 1535
rect 3189 1481 3213 1515
rect 3247 1481 3261 1515
rect 3189 1315 3261 1481
rect 3535 1515 3607 1535
rect 3535 1481 3549 1515
rect 3583 1481 3607 1515
rect 3189 1281 3213 1315
rect 3247 1281 3261 1315
rect 3189 1261 3261 1281
rect 3535 1315 3607 1481
rect 3535 1281 3549 1315
rect 3583 1281 3607 1315
rect 3535 1261 3607 1281
rect 3189 1247 3607 1261
rect 3189 1213 3213 1247
rect 3247 1213 3281 1247
rect 3315 1213 3481 1247
rect 3515 1213 3549 1247
rect 3583 1213 3607 1247
rect 3189 1189 3607 1213
rect -3811 583 -3393 607
rect -3811 549 -3787 583
rect -3753 549 -3719 583
rect -3685 549 -3519 583
rect -3485 549 -3451 583
rect -3417 549 -3393 583
rect -3811 535 -3393 549
rect -3811 515 -3739 535
rect -3811 481 -3787 515
rect -3753 481 -3739 515
rect -3811 315 -3739 481
rect -3465 515 -3393 535
rect -3465 481 -3451 515
rect -3417 481 -3393 515
rect -3811 281 -3787 315
rect -3753 281 -3739 315
rect -3811 261 -3739 281
rect -3465 315 -3393 481
rect -3465 281 -3451 315
rect -3417 281 -3393 315
rect -3465 261 -3393 281
rect -3811 247 -3393 261
rect -3811 213 -3787 247
rect -3753 213 -3719 247
rect -3685 213 -3519 247
rect -3485 213 -3451 247
rect -3417 213 -3393 247
rect -3811 189 -3393 213
rect -2811 583 -2393 607
rect -2811 549 -2787 583
rect -2753 549 -2719 583
rect -2685 549 -2519 583
rect -2485 549 -2451 583
rect -2417 549 -2393 583
rect -2811 535 -2393 549
rect -2811 515 -2739 535
rect -2811 481 -2787 515
rect -2753 481 -2739 515
rect -2811 315 -2739 481
rect -2465 515 -2393 535
rect -2465 481 -2451 515
rect -2417 481 -2393 515
rect -2811 281 -2787 315
rect -2753 281 -2739 315
rect -2811 261 -2739 281
rect -2465 315 -2393 481
rect -2465 281 -2451 315
rect -2417 281 -2393 315
rect -2465 261 -2393 281
rect -2811 247 -2393 261
rect -2811 213 -2787 247
rect -2753 213 -2719 247
rect -2685 213 -2519 247
rect -2485 213 -2451 247
rect -2417 213 -2393 247
rect -2811 189 -2393 213
rect -1811 583 -1393 607
rect -1811 549 -1787 583
rect -1753 549 -1719 583
rect -1685 549 -1519 583
rect -1485 549 -1451 583
rect -1417 549 -1393 583
rect -1811 535 -1393 549
rect -1811 515 -1739 535
rect -1811 481 -1787 515
rect -1753 481 -1739 515
rect -1811 315 -1739 481
rect -1465 515 -1393 535
rect -1465 481 -1451 515
rect -1417 481 -1393 515
rect -1811 281 -1787 315
rect -1753 281 -1739 315
rect -1811 261 -1739 281
rect -1465 315 -1393 481
rect -1465 281 -1451 315
rect -1417 281 -1393 315
rect -1465 261 -1393 281
rect -1811 247 -1393 261
rect -1811 213 -1787 247
rect -1753 213 -1719 247
rect -1685 213 -1519 247
rect -1485 213 -1451 247
rect -1417 213 -1393 247
rect -1811 189 -1393 213
rect -811 583 -393 607
rect -811 549 -787 583
rect -753 549 -719 583
rect -685 549 -519 583
rect -485 549 -451 583
rect -417 549 -393 583
rect -811 535 -393 549
rect -811 515 -739 535
rect -811 481 -787 515
rect -753 481 -739 515
rect -811 315 -739 481
rect -465 515 -393 535
rect -465 481 -451 515
rect -417 481 -393 515
rect -811 281 -787 315
rect -753 281 -739 315
rect -811 261 -739 281
rect -465 315 -393 481
rect -465 281 -451 315
rect -417 281 -393 315
rect -465 261 -393 281
rect -811 247 -393 261
rect -811 213 -787 247
rect -753 213 -719 247
rect -685 213 -519 247
rect -485 213 -451 247
rect -417 213 -393 247
rect -811 189 -393 213
rect 1189 583 1607 607
rect 1189 549 1213 583
rect 1247 549 1281 583
rect 1315 549 1481 583
rect 1515 549 1549 583
rect 1583 549 1607 583
rect 1189 535 1607 549
rect 1189 515 1261 535
rect 1189 481 1213 515
rect 1247 481 1261 515
rect 1189 315 1261 481
rect 1535 515 1607 535
rect 1535 481 1549 515
rect 1583 481 1607 515
rect 1189 281 1213 315
rect 1247 281 1261 315
rect 1189 261 1261 281
rect 1535 315 1607 481
rect 1535 281 1549 315
rect 1583 281 1607 315
rect 1535 261 1607 281
rect 1189 247 1607 261
rect 1189 213 1213 247
rect 1247 213 1281 247
rect 1315 213 1481 247
rect 1515 213 1549 247
rect 1583 213 1607 247
rect 1189 189 1607 213
rect 2189 583 2607 607
rect 2189 549 2213 583
rect 2247 549 2281 583
rect 2315 549 2481 583
rect 2515 549 2549 583
rect 2583 549 2607 583
rect 2189 535 2607 549
rect 2189 515 2261 535
rect 2189 481 2213 515
rect 2247 481 2261 515
rect 2189 315 2261 481
rect 2535 515 2607 535
rect 2535 481 2549 515
rect 2583 481 2607 515
rect 2189 281 2213 315
rect 2247 281 2261 315
rect 2189 261 2261 281
rect 2535 315 2607 481
rect 2535 281 2549 315
rect 2583 281 2607 315
rect 2535 261 2607 281
rect 2189 247 2607 261
rect 2189 213 2213 247
rect 2247 213 2281 247
rect 2315 213 2481 247
rect 2515 213 2549 247
rect 2583 213 2607 247
rect 2189 189 2607 213
rect 3189 583 3607 607
rect 3189 549 3213 583
rect 3247 549 3281 583
rect 3315 549 3481 583
rect 3515 549 3549 583
rect 3583 549 3607 583
rect 3189 535 3607 549
rect 3189 515 3261 535
rect 3189 481 3213 515
rect 3247 481 3261 515
rect 3189 315 3261 481
rect 3535 515 3607 535
rect 3535 481 3549 515
rect 3583 481 3607 515
rect 3189 281 3213 315
rect 3247 281 3261 315
rect 3189 261 3261 281
rect 3535 315 3607 481
rect 3535 281 3549 315
rect 3583 281 3607 315
rect 3535 261 3607 281
rect 3189 247 3607 261
rect 3189 213 3213 247
rect 3247 213 3281 247
rect 3315 213 3481 247
rect 3515 213 3549 247
rect 3583 213 3607 247
rect 3189 189 3607 213
rect -3811 -417 -3393 -393
rect -3811 -451 -3787 -417
rect -3753 -451 -3719 -417
rect -3685 -451 -3519 -417
rect -3485 -451 -3451 -417
rect -3417 -451 -3393 -417
rect -3811 -465 -3393 -451
rect -3811 -485 -3739 -465
rect -3811 -519 -3787 -485
rect -3753 -519 -3739 -485
rect -3811 -685 -3739 -519
rect -3465 -485 -3393 -465
rect -3465 -519 -3451 -485
rect -3417 -519 -3393 -485
rect -3811 -719 -3787 -685
rect -3753 -719 -3739 -685
rect -3811 -739 -3739 -719
rect -3465 -685 -3393 -519
rect -3465 -719 -3451 -685
rect -3417 -719 -3393 -685
rect -3465 -739 -3393 -719
rect -3811 -753 -3393 -739
rect -3811 -787 -3787 -753
rect -3753 -787 -3719 -753
rect -3685 -787 -3519 -753
rect -3485 -787 -3451 -753
rect -3417 -787 -3393 -753
rect -3811 -811 -3393 -787
rect -2811 -417 -2393 -393
rect -2811 -451 -2787 -417
rect -2753 -451 -2719 -417
rect -2685 -451 -2519 -417
rect -2485 -451 -2451 -417
rect -2417 -451 -2393 -417
rect -2811 -465 -2393 -451
rect -2811 -485 -2739 -465
rect -2811 -519 -2787 -485
rect -2753 -519 -2739 -485
rect -2811 -685 -2739 -519
rect -2465 -485 -2393 -465
rect -2465 -519 -2451 -485
rect -2417 -519 -2393 -485
rect -2811 -719 -2787 -685
rect -2753 -719 -2739 -685
rect -2811 -739 -2739 -719
rect -2465 -685 -2393 -519
rect -2465 -719 -2451 -685
rect -2417 -719 -2393 -685
rect -2465 -739 -2393 -719
rect -2811 -753 -2393 -739
rect -2811 -787 -2787 -753
rect -2753 -787 -2719 -753
rect -2685 -787 -2519 -753
rect -2485 -787 -2451 -753
rect -2417 -787 -2393 -753
rect -2811 -811 -2393 -787
rect -1811 -417 -1393 -393
rect -1811 -451 -1787 -417
rect -1753 -451 -1719 -417
rect -1685 -451 -1519 -417
rect -1485 -451 -1451 -417
rect -1417 -451 -1393 -417
rect -1811 -465 -1393 -451
rect -1811 -485 -1739 -465
rect -1811 -519 -1787 -485
rect -1753 -519 -1739 -485
rect -1811 -685 -1739 -519
rect -1465 -485 -1393 -465
rect -1465 -519 -1451 -485
rect -1417 -519 -1393 -485
rect -1811 -719 -1787 -685
rect -1753 -719 -1739 -685
rect -1811 -739 -1739 -719
rect -1465 -685 -1393 -519
rect -1465 -719 -1451 -685
rect -1417 -719 -1393 -685
rect -1465 -739 -1393 -719
rect -1811 -753 -1393 -739
rect -1811 -787 -1787 -753
rect -1753 -787 -1719 -753
rect -1685 -787 -1519 -753
rect -1485 -787 -1451 -753
rect -1417 -787 -1393 -753
rect -1811 -811 -1393 -787
rect -811 -417 -393 -393
rect -811 -451 -787 -417
rect -753 -451 -719 -417
rect -685 -451 -519 -417
rect -485 -451 -451 -417
rect -417 -451 -393 -417
rect -811 -465 -393 -451
rect -811 -485 -739 -465
rect -811 -519 -787 -485
rect -753 -519 -739 -485
rect -811 -685 -739 -519
rect -465 -485 -393 -465
rect -465 -519 -451 -485
rect -417 -519 -393 -485
rect -811 -719 -787 -685
rect -753 -719 -739 -685
rect -811 -739 -739 -719
rect -465 -685 -393 -519
rect -465 -719 -451 -685
rect -417 -719 -393 -685
rect -465 -739 -393 -719
rect -811 -753 -393 -739
rect -811 -787 -787 -753
rect -753 -787 -719 -753
rect -685 -787 -519 -753
rect -485 -787 -451 -753
rect -417 -787 -393 -753
rect -811 -811 -393 -787
rect 189 -417 607 -393
rect 189 -451 213 -417
rect 247 -451 281 -417
rect 315 -451 481 -417
rect 515 -451 549 -417
rect 583 -451 607 -417
rect 189 -465 607 -451
rect 189 -485 261 -465
rect 189 -519 213 -485
rect 247 -519 261 -485
rect 189 -685 261 -519
rect 535 -485 607 -465
rect 535 -519 549 -485
rect 583 -519 607 -485
rect 189 -719 213 -685
rect 247 -719 261 -685
rect 189 -739 261 -719
rect 535 -685 607 -519
rect 535 -719 549 -685
rect 583 -719 607 -685
rect 535 -739 607 -719
rect 189 -753 607 -739
rect 189 -787 213 -753
rect 247 -787 281 -753
rect 315 -787 481 -753
rect 515 -787 549 -753
rect 583 -787 607 -753
rect 189 -811 607 -787
rect 1189 -417 1607 -393
rect 1189 -451 1213 -417
rect 1247 -451 1281 -417
rect 1315 -451 1481 -417
rect 1515 -451 1549 -417
rect 1583 -451 1607 -417
rect 1189 -465 1607 -451
rect 1189 -485 1261 -465
rect 1189 -519 1213 -485
rect 1247 -519 1261 -485
rect 1189 -685 1261 -519
rect 1535 -485 1607 -465
rect 1535 -519 1549 -485
rect 1583 -519 1607 -485
rect 1189 -719 1213 -685
rect 1247 -719 1261 -685
rect 1189 -739 1261 -719
rect 1535 -685 1607 -519
rect 1535 -719 1549 -685
rect 1583 -719 1607 -685
rect 1535 -739 1607 -719
rect 1189 -753 1607 -739
rect 1189 -787 1213 -753
rect 1247 -787 1281 -753
rect 1315 -787 1481 -753
rect 1515 -787 1549 -753
rect 1583 -787 1607 -753
rect 1189 -811 1607 -787
rect 2189 -417 2607 -393
rect 2189 -451 2213 -417
rect 2247 -451 2281 -417
rect 2315 -451 2481 -417
rect 2515 -451 2549 -417
rect 2583 -451 2607 -417
rect 2189 -465 2607 -451
rect 2189 -485 2261 -465
rect 2189 -519 2213 -485
rect 2247 -519 2261 -485
rect 2189 -685 2261 -519
rect 2535 -485 2607 -465
rect 2535 -519 2549 -485
rect 2583 -519 2607 -485
rect 2189 -719 2213 -685
rect 2247 -719 2261 -685
rect 2189 -739 2261 -719
rect 2535 -685 2607 -519
rect 2535 -719 2549 -685
rect 2583 -719 2607 -685
rect 2535 -739 2607 -719
rect 2189 -753 2607 -739
rect 2189 -787 2213 -753
rect 2247 -787 2281 -753
rect 2315 -787 2481 -753
rect 2515 -787 2549 -753
rect 2583 -787 2607 -753
rect 2189 -811 2607 -787
rect 3189 -417 3607 -393
rect 3189 -451 3213 -417
rect 3247 -451 3281 -417
rect 3315 -451 3481 -417
rect 3515 -451 3549 -417
rect 3583 -451 3607 -417
rect 3189 -465 3607 -451
rect 3189 -485 3261 -465
rect 3189 -519 3213 -485
rect 3247 -519 3261 -485
rect 3189 -685 3261 -519
rect 3535 -485 3607 -465
rect 3535 -519 3549 -485
rect 3583 -519 3607 -485
rect 3189 -719 3213 -685
rect 3247 -719 3261 -685
rect 3189 -739 3261 -719
rect 3535 -685 3607 -519
rect 3535 -719 3549 -685
rect 3583 -719 3607 -685
rect 3535 -739 3607 -719
rect 3189 -753 3607 -739
rect 3189 -787 3213 -753
rect 3247 -787 3281 -753
rect 3315 -787 3481 -753
rect 3515 -787 3549 -753
rect 3583 -787 3607 -753
rect 3189 -811 3607 -787
rect -811 -1417 -393 -1393
rect -811 -1451 -787 -1417
rect -753 -1451 -719 -1417
rect -685 -1451 -519 -1417
rect -485 -1451 -451 -1417
rect -417 -1451 -393 -1417
rect -811 -1465 -393 -1451
rect -811 -1485 -739 -1465
rect -811 -1519 -787 -1485
rect -753 -1519 -739 -1485
rect -811 -1685 -739 -1519
rect -465 -1485 -393 -1465
rect -465 -1519 -451 -1485
rect -417 -1519 -393 -1485
rect -811 -1719 -787 -1685
rect -753 -1719 -739 -1685
rect -811 -1739 -739 -1719
rect -465 -1685 -393 -1519
rect -465 -1719 -451 -1685
rect -417 -1719 -393 -1685
rect -465 -1739 -393 -1719
rect -811 -1753 -393 -1739
rect -811 -1787 -787 -1753
rect -753 -1787 -719 -1753
rect -685 -1787 -519 -1753
rect -485 -1787 -451 -1753
rect -417 -1787 -393 -1753
rect -811 -1811 -393 -1787
rect 189 -1417 607 -1393
rect 189 -1451 213 -1417
rect 247 -1451 281 -1417
rect 315 -1451 481 -1417
rect 515 -1451 549 -1417
rect 583 -1451 607 -1417
rect 189 -1465 607 -1451
rect 189 -1485 261 -1465
rect 189 -1519 213 -1485
rect 247 -1519 261 -1485
rect 189 -1685 261 -1519
rect 535 -1485 607 -1465
rect 535 -1519 549 -1485
rect 583 -1519 607 -1485
rect 189 -1719 213 -1685
rect 247 -1719 261 -1685
rect 189 -1739 261 -1719
rect 535 -1685 607 -1519
rect 535 -1719 549 -1685
rect 583 -1719 607 -1685
rect 535 -1739 607 -1719
rect 189 -1753 607 -1739
rect 189 -1787 213 -1753
rect 247 -1787 281 -1753
rect 315 -1787 481 -1753
rect 515 -1787 549 -1753
rect 583 -1787 607 -1753
rect 189 -1811 607 -1787
rect 1189 -1417 1607 -1393
rect 1189 -1451 1213 -1417
rect 1247 -1451 1281 -1417
rect 1315 -1451 1481 -1417
rect 1515 -1451 1549 -1417
rect 1583 -1451 1607 -1417
rect 1189 -1465 1607 -1451
rect 1189 -1485 1261 -1465
rect 1189 -1519 1213 -1485
rect 1247 -1519 1261 -1485
rect 1189 -1685 1261 -1519
rect 1535 -1485 1607 -1465
rect 1535 -1519 1549 -1485
rect 1583 -1519 1607 -1485
rect 1189 -1719 1213 -1685
rect 1247 -1719 1261 -1685
rect 1189 -1739 1261 -1719
rect 1535 -1685 1607 -1519
rect 1535 -1719 1549 -1685
rect 1583 -1719 1607 -1685
rect 1535 -1739 1607 -1719
rect 1189 -1753 1607 -1739
rect 1189 -1787 1213 -1753
rect 1247 -1787 1281 -1753
rect 1315 -1787 1481 -1753
rect 1515 -1787 1549 -1753
rect 1583 -1787 1607 -1753
rect 1189 -1811 1607 -1787
rect 2189 -1417 2607 -1393
rect 2189 -1451 2213 -1417
rect 2247 -1451 2281 -1417
rect 2315 -1451 2481 -1417
rect 2515 -1451 2549 -1417
rect 2583 -1451 2607 -1417
rect 2189 -1465 2607 -1451
rect 2189 -1485 2261 -1465
rect 2189 -1519 2213 -1485
rect 2247 -1519 2261 -1485
rect 2189 -1685 2261 -1519
rect 2535 -1485 2607 -1465
rect 2535 -1519 2549 -1485
rect 2583 -1519 2607 -1485
rect 2189 -1719 2213 -1685
rect 2247 -1719 2261 -1685
rect 2189 -1739 2261 -1719
rect 2535 -1685 2607 -1519
rect 2535 -1719 2549 -1685
rect 2583 -1719 2607 -1685
rect 2535 -1739 2607 -1719
rect 2189 -1753 2607 -1739
rect 2189 -1787 2213 -1753
rect 2247 -1787 2281 -1753
rect 2315 -1787 2481 -1753
rect 2515 -1787 2549 -1753
rect 2583 -1787 2607 -1753
rect 2189 -1811 2607 -1787
rect 3189 -1417 3607 -1393
rect 3189 -1451 3213 -1417
rect 3247 -1451 3281 -1417
rect 3315 -1451 3481 -1417
rect 3515 -1451 3549 -1417
rect 3583 -1451 3607 -1417
rect 3189 -1465 3607 -1451
rect 3189 -1485 3261 -1465
rect 3189 -1519 3213 -1485
rect 3247 -1519 3261 -1485
rect 3189 -1685 3261 -1519
rect 3535 -1485 3607 -1465
rect 3535 -1519 3549 -1485
rect 3583 -1519 3607 -1485
rect 3189 -1719 3213 -1685
rect 3247 -1719 3261 -1685
rect 3189 -1739 3261 -1719
rect 3535 -1685 3607 -1519
rect 3535 -1719 3549 -1685
rect 3583 -1719 3607 -1685
rect 3535 -1739 3607 -1719
rect 3189 -1753 3607 -1739
rect 3189 -1787 3213 -1753
rect 3247 -1787 3281 -1753
rect 3315 -1787 3481 -1753
rect 3515 -1787 3549 -1753
rect 3583 -1787 3607 -1753
rect 3189 -1811 3607 -1787
rect -811 -2417 -393 -2393
rect -811 -2451 -787 -2417
rect -753 -2451 -719 -2417
rect -685 -2451 -519 -2417
rect -485 -2451 -451 -2417
rect -417 -2451 -393 -2417
rect -811 -2465 -393 -2451
rect -811 -2485 -739 -2465
rect -811 -2519 -787 -2485
rect -753 -2519 -739 -2485
rect -811 -2685 -739 -2519
rect -465 -2485 -393 -2465
rect -465 -2519 -451 -2485
rect -417 -2519 -393 -2485
rect -811 -2719 -787 -2685
rect -753 -2719 -739 -2685
rect -811 -2739 -739 -2719
rect -465 -2685 -393 -2519
rect -465 -2719 -451 -2685
rect -417 -2719 -393 -2685
rect -465 -2739 -393 -2719
rect -811 -2753 -393 -2739
rect -811 -2787 -787 -2753
rect -753 -2787 -719 -2753
rect -685 -2787 -519 -2753
rect -485 -2787 -451 -2753
rect -417 -2787 -393 -2753
rect -811 -2811 -393 -2787
rect 189 -2417 607 -2393
rect 189 -2451 213 -2417
rect 247 -2451 281 -2417
rect 315 -2451 481 -2417
rect 515 -2451 549 -2417
rect 583 -2451 607 -2417
rect 189 -2465 607 -2451
rect 189 -2485 261 -2465
rect 189 -2519 213 -2485
rect 247 -2519 261 -2485
rect 189 -2685 261 -2519
rect 535 -2485 607 -2465
rect 535 -2519 549 -2485
rect 583 -2519 607 -2485
rect 189 -2719 213 -2685
rect 247 -2719 261 -2685
rect 189 -2739 261 -2719
rect 535 -2685 607 -2519
rect 535 -2719 549 -2685
rect 583 -2719 607 -2685
rect 535 -2739 607 -2719
rect 189 -2753 607 -2739
rect 189 -2787 213 -2753
rect 247 -2787 281 -2753
rect 315 -2787 481 -2753
rect 515 -2787 549 -2753
rect 583 -2787 607 -2753
rect 189 -2811 607 -2787
rect 1189 -2417 1607 -2393
rect 1189 -2451 1213 -2417
rect 1247 -2451 1281 -2417
rect 1315 -2451 1481 -2417
rect 1515 -2451 1549 -2417
rect 1583 -2451 1607 -2417
rect 1189 -2465 1607 -2451
rect 1189 -2485 1261 -2465
rect 1189 -2519 1213 -2485
rect 1247 -2519 1261 -2485
rect 1189 -2685 1261 -2519
rect 1535 -2485 1607 -2465
rect 1535 -2519 1549 -2485
rect 1583 -2519 1607 -2485
rect 1189 -2719 1213 -2685
rect 1247 -2719 1261 -2685
rect 1189 -2739 1261 -2719
rect 1535 -2685 1607 -2519
rect 1535 -2719 1549 -2685
rect 1583 -2719 1607 -2685
rect 1535 -2739 1607 -2719
rect 1189 -2753 1607 -2739
rect 1189 -2787 1213 -2753
rect 1247 -2787 1281 -2753
rect 1315 -2787 1481 -2753
rect 1515 -2787 1549 -2753
rect 1583 -2787 1607 -2753
rect 1189 -2811 1607 -2787
rect 2189 -2417 2607 -2393
rect 2189 -2451 2213 -2417
rect 2247 -2451 2281 -2417
rect 2315 -2451 2481 -2417
rect 2515 -2451 2549 -2417
rect 2583 -2451 2607 -2417
rect 2189 -2465 2607 -2451
rect 2189 -2485 2261 -2465
rect 2189 -2519 2213 -2485
rect 2247 -2519 2261 -2485
rect 2189 -2685 2261 -2519
rect 2535 -2485 2607 -2465
rect 2535 -2519 2549 -2485
rect 2583 -2519 2607 -2485
rect 2189 -2719 2213 -2685
rect 2247 -2719 2261 -2685
rect 2189 -2739 2261 -2719
rect 2535 -2685 2607 -2519
rect 2535 -2719 2549 -2685
rect 2583 -2719 2607 -2685
rect 2535 -2739 2607 -2719
rect 2189 -2753 2607 -2739
rect 2189 -2787 2213 -2753
rect 2247 -2787 2281 -2753
rect 2315 -2787 2481 -2753
rect 2515 -2787 2549 -2753
rect 2583 -2787 2607 -2753
rect 2189 -2811 2607 -2787
rect 3189 -2417 3607 -2393
rect 3189 -2451 3213 -2417
rect 3247 -2451 3281 -2417
rect 3315 -2451 3481 -2417
rect 3515 -2451 3549 -2417
rect 3583 -2451 3607 -2417
rect 3189 -2465 3607 -2451
rect 3189 -2485 3261 -2465
rect 3189 -2519 3213 -2485
rect 3247 -2519 3261 -2485
rect 3189 -2685 3261 -2519
rect 3535 -2485 3607 -2465
rect 3535 -2519 3549 -2485
rect 3583 -2519 3607 -2485
rect 3189 -2719 3213 -2685
rect 3247 -2719 3261 -2685
rect 3189 -2739 3261 -2719
rect 3535 -2685 3607 -2519
rect 3535 -2719 3549 -2685
rect 3583 -2719 3607 -2685
rect 3535 -2739 3607 -2719
rect 3189 -2753 3607 -2739
rect 3189 -2787 3213 -2753
rect 3247 -2787 3281 -2753
rect 3315 -2787 3481 -2753
rect 3515 -2787 3549 -2753
rect 3583 -2787 3607 -2753
rect 3189 -2811 3607 -2787
<< psubdiffcont >>
rect -3940 1702 -3906 1736
rect -3872 1702 -3838 1736
rect -3804 1702 -3770 1736
rect -3736 1702 -3702 1736
rect -3502 1702 -3468 1736
rect -3434 1702 -3400 1736
rect -3366 1702 -3332 1736
rect -3298 1702 -3264 1736
rect -3940 1634 -3906 1668
rect -3298 1634 -3264 1668
rect -3940 1566 -3906 1600
rect -3940 1498 -3906 1532
rect -3940 1264 -3906 1298
rect -3940 1196 -3906 1230
rect -3298 1566 -3264 1600
rect -3298 1498 -3264 1532
rect -3298 1264 -3264 1298
rect -3298 1196 -3264 1230
rect -3940 1128 -3906 1162
rect -3298 1128 -3264 1162
rect -3940 1060 -3906 1094
rect -3872 1060 -3838 1094
rect -3804 1060 -3770 1094
rect -3736 1060 -3702 1094
rect -3502 1060 -3468 1094
rect -3434 1060 -3400 1094
rect -3366 1060 -3332 1094
rect -3298 1060 -3264 1094
rect -2940 1702 -2906 1736
rect -2872 1702 -2838 1736
rect -2804 1702 -2770 1736
rect -2736 1702 -2702 1736
rect -2502 1702 -2468 1736
rect -2434 1702 -2400 1736
rect -2366 1702 -2332 1736
rect -2298 1702 -2264 1736
rect -2940 1634 -2906 1668
rect -2298 1634 -2264 1668
rect -2940 1566 -2906 1600
rect -2940 1498 -2906 1532
rect -2940 1264 -2906 1298
rect -2940 1196 -2906 1230
rect -2298 1566 -2264 1600
rect -2298 1498 -2264 1532
rect -2298 1264 -2264 1298
rect -2298 1196 -2264 1230
rect -2940 1128 -2906 1162
rect -2298 1128 -2264 1162
rect -2940 1060 -2906 1094
rect -2872 1060 -2838 1094
rect -2804 1060 -2770 1094
rect -2736 1060 -2702 1094
rect -2502 1060 -2468 1094
rect -2434 1060 -2400 1094
rect -2366 1060 -2332 1094
rect -2298 1060 -2264 1094
rect -1940 1702 -1906 1736
rect -1872 1702 -1838 1736
rect -1804 1702 -1770 1736
rect -1736 1702 -1702 1736
rect -1502 1702 -1468 1736
rect -1434 1702 -1400 1736
rect -1366 1702 -1332 1736
rect -1298 1702 -1264 1736
rect -1940 1634 -1906 1668
rect -1298 1634 -1264 1668
rect -1940 1566 -1906 1600
rect -1940 1498 -1906 1532
rect -1940 1264 -1906 1298
rect -1940 1196 -1906 1230
rect -1298 1566 -1264 1600
rect -1298 1498 -1264 1532
rect -1298 1264 -1264 1298
rect -1298 1196 -1264 1230
rect -1940 1128 -1906 1162
rect -1298 1128 -1264 1162
rect -1940 1060 -1906 1094
rect -1872 1060 -1838 1094
rect -1804 1060 -1770 1094
rect -1736 1060 -1702 1094
rect -1502 1060 -1468 1094
rect -1434 1060 -1400 1094
rect -1366 1060 -1332 1094
rect -1298 1060 -1264 1094
rect -940 1702 -906 1736
rect -872 1702 -838 1736
rect -804 1702 -770 1736
rect -736 1702 -702 1736
rect -502 1702 -468 1736
rect -434 1702 -400 1736
rect -366 1702 -332 1736
rect -298 1702 -264 1736
rect -940 1634 -906 1668
rect -298 1634 -264 1668
rect -940 1566 -906 1600
rect -940 1498 -906 1532
rect -940 1264 -906 1298
rect -940 1196 -906 1230
rect -298 1566 -264 1600
rect -298 1498 -264 1532
rect -298 1264 -264 1298
rect -298 1196 -264 1230
rect -940 1128 -906 1162
rect -298 1128 -264 1162
rect -940 1060 -906 1094
rect -872 1060 -838 1094
rect -804 1060 -770 1094
rect -736 1060 -702 1094
rect -502 1060 -468 1094
rect -434 1060 -400 1094
rect -366 1060 -332 1094
rect -298 1060 -264 1094
rect 60 1702 94 1736
rect 128 1702 162 1736
rect 196 1702 230 1736
rect 264 1702 298 1736
rect 498 1702 532 1736
rect 566 1702 600 1736
rect 634 1702 668 1736
rect 702 1702 736 1736
rect 60 1634 94 1668
rect 702 1634 736 1668
rect 60 1566 94 1600
rect 60 1498 94 1532
rect 60 1264 94 1298
rect 60 1196 94 1230
rect 702 1566 736 1600
rect 702 1498 736 1532
rect 702 1264 736 1298
rect 702 1196 736 1230
rect 60 1128 94 1162
rect 702 1128 736 1162
rect 60 1060 94 1094
rect 128 1060 162 1094
rect 196 1060 230 1094
rect 264 1060 298 1094
rect 498 1060 532 1094
rect 566 1060 600 1094
rect 634 1060 668 1094
rect 702 1060 736 1094
rect 1060 1702 1094 1736
rect 1128 1702 1162 1736
rect 1196 1702 1230 1736
rect 1264 1702 1298 1736
rect 1498 1702 1532 1736
rect 1566 1702 1600 1736
rect 1634 1702 1668 1736
rect 1702 1702 1736 1736
rect 1060 1634 1094 1668
rect 1702 1634 1736 1668
rect 1060 1566 1094 1600
rect 1060 1498 1094 1532
rect 1060 1264 1094 1298
rect 1060 1196 1094 1230
rect 1702 1566 1736 1600
rect 1702 1498 1736 1532
rect 1702 1264 1736 1298
rect 1702 1196 1736 1230
rect 1060 1128 1094 1162
rect 1702 1128 1736 1162
rect 1060 1060 1094 1094
rect 1128 1060 1162 1094
rect 1196 1060 1230 1094
rect 1264 1060 1298 1094
rect 1498 1060 1532 1094
rect 1566 1060 1600 1094
rect 1634 1060 1668 1094
rect 1702 1060 1736 1094
rect 2060 1702 2094 1736
rect 2128 1702 2162 1736
rect 2196 1702 2230 1736
rect 2264 1702 2298 1736
rect 2498 1702 2532 1736
rect 2566 1702 2600 1736
rect 2634 1702 2668 1736
rect 2702 1702 2736 1736
rect 2060 1634 2094 1668
rect 2702 1634 2736 1668
rect 2060 1566 2094 1600
rect 2060 1498 2094 1532
rect 2060 1264 2094 1298
rect 2060 1196 2094 1230
rect 2702 1566 2736 1600
rect 2702 1498 2736 1532
rect 2702 1264 2736 1298
rect 2702 1196 2736 1230
rect 2060 1128 2094 1162
rect 2702 1128 2736 1162
rect 2060 1060 2094 1094
rect 2128 1060 2162 1094
rect 2196 1060 2230 1094
rect 2264 1060 2298 1094
rect 2498 1060 2532 1094
rect 2566 1060 2600 1094
rect 2634 1060 2668 1094
rect 2702 1060 2736 1094
rect 3060 1702 3094 1736
rect 3128 1702 3162 1736
rect 3196 1702 3230 1736
rect 3264 1702 3298 1736
rect 3498 1702 3532 1736
rect 3566 1702 3600 1736
rect 3634 1702 3668 1736
rect 3702 1702 3736 1736
rect 3060 1634 3094 1668
rect 3702 1634 3736 1668
rect 3060 1566 3094 1600
rect 3060 1498 3094 1532
rect 3060 1264 3094 1298
rect 3060 1196 3094 1230
rect 3702 1566 3736 1600
rect 3702 1498 3736 1532
rect 3702 1264 3736 1298
rect 3702 1196 3736 1230
rect 3060 1128 3094 1162
rect 3702 1128 3736 1162
rect 3060 1060 3094 1094
rect 3128 1060 3162 1094
rect 3196 1060 3230 1094
rect 3264 1060 3298 1094
rect 3498 1060 3532 1094
rect 3566 1060 3600 1094
rect 3634 1060 3668 1094
rect 3702 1060 3736 1094
rect -3940 702 -3906 736
rect -3872 702 -3838 736
rect -3804 702 -3770 736
rect -3736 702 -3702 736
rect -3502 702 -3468 736
rect -3434 702 -3400 736
rect -3366 702 -3332 736
rect -3298 702 -3264 736
rect -3940 634 -3906 668
rect -3298 634 -3264 668
rect -3940 566 -3906 600
rect -3940 498 -3906 532
rect -3940 264 -3906 298
rect -3940 196 -3906 230
rect -3298 566 -3264 600
rect -3298 498 -3264 532
rect -3298 264 -3264 298
rect -3298 196 -3264 230
rect -3940 128 -3906 162
rect -3298 128 -3264 162
rect -3940 60 -3906 94
rect -3872 60 -3838 94
rect -3804 60 -3770 94
rect -3736 60 -3702 94
rect -3502 60 -3468 94
rect -3434 60 -3400 94
rect -3366 60 -3332 94
rect -3298 60 -3264 94
rect -2940 702 -2906 736
rect -2872 702 -2838 736
rect -2804 702 -2770 736
rect -2736 702 -2702 736
rect -2502 702 -2468 736
rect -2434 702 -2400 736
rect -2366 702 -2332 736
rect -2298 702 -2264 736
rect -2940 634 -2906 668
rect -2298 634 -2264 668
rect -2940 566 -2906 600
rect -2940 498 -2906 532
rect -2940 264 -2906 298
rect -2940 196 -2906 230
rect -2298 566 -2264 600
rect -2298 498 -2264 532
rect -2298 264 -2264 298
rect -2298 196 -2264 230
rect -2940 128 -2906 162
rect -2298 128 -2264 162
rect -2940 60 -2906 94
rect -2872 60 -2838 94
rect -2804 60 -2770 94
rect -2736 60 -2702 94
rect -2502 60 -2468 94
rect -2434 60 -2400 94
rect -2366 60 -2332 94
rect -2298 60 -2264 94
rect -1940 702 -1906 736
rect -1872 702 -1838 736
rect -1804 702 -1770 736
rect -1736 702 -1702 736
rect -1502 702 -1468 736
rect -1434 702 -1400 736
rect -1366 702 -1332 736
rect -1298 702 -1264 736
rect -1940 634 -1906 668
rect -1298 634 -1264 668
rect -1940 566 -1906 600
rect -1940 498 -1906 532
rect -1940 264 -1906 298
rect -1940 196 -1906 230
rect -1298 566 -1264 600
rect -1298 498 -1264 532
rect -1298 264 -1264 298
rect -1298 196 -1264 230
rect -1940 128 -1906 162
rect -1298 128 -1264 162
rect -1940 60 -1906 94
rect -1872 60 -1838 94
rect -1804 60 -1770 94
rect -1736 60 -1702 94
rect -1502 60 -1468 94
rect -1434 60 -1400 94
rect -1366 60 -1332 94
rect -1298 60 -1264 94
rect -940 702 -906 736
rect -872 702 -838 736
rect -804 702 -770 736
rect -736 702 -702 736
rect -502 702 -468 736
rect -434 702 -400 736
rect -366 702 -332 736
rect -298 702 -264 736
rect -940 634 -906 668
rect -298 634 -264 668
rect -940 566 -906 600
rect -940 498 -906 532
rect -940 264 -906 298
rect -940 196 -906 230
rect -298 566 -264 600
rect -298 498 -264 532
rect -298 264 -264 298
rect -298 196 -264 230
rect -940 128 -906 162
rect -298 128 -264 162
rect -940 60 -906 94
rect -872 60 -838 94
rect -804 60 -770 94
rect -736 60 -702 94
rect -502 60 -468 94
rect -434 60 -400 94
rect -366 60 -332 94
rect -298 60 -264 94
rect 1060 702 1094 736
rect 1128 702 1162 736
rect 1196 702 1230 736
rect 1264 702 1298 736
rect 1498 702 1532 736
rect 1566 702 1600 736
rect 1634 702 1668 736
rect 1702 702 1736 736
rect 1060 634 1094 668
rect 1702 634 1736 668
rect 1060 566 1094 600
rect 1060 498 1094 532
rect 1060 264 1094 298
rect 1060 196 1094 230
rect 1702 566 1736 600
rect 1702 498 1736 532
rect 1702 264 1736 298
rect 1702 196 1736 230
rect 1060 128 1094 162
rect 1702 128 1736 162
rect 1060 60 1094 94
rect 1128 60 1162 94
rect 1196 60 1230 94
rect 1264 60 1298 94
rect 1498 60 1532 94
rect 1566 60 1600 94
rect 1634 60 1668 94
rect 1702 60 1736 94
rect 2060 702 2094 736
rect 2128 702 2162 736
rect 2196 702 2230 736
rect 2264 702 2298 736
rect 2498 702 2532 736
rect 2566 702 2600 736
rect 2634 702 2668 736
rect 2702 702 2736 736
rect 2060 634 2094 668
rect 2702 634 2736 668
rect 2060 566 2094 600
rect 2060 498 2094 532
rect 2060 264 2094 298
rect 2060 196 2094 230
rect 2702 566 2736 600
rect 2702 498 2736 532
rect 2702 264 2736 298
rect 2702 196 2736 230
rect 2060 128 2094 162
rect 2702 128 2736 162
rect 2060 60 2094 94
rect 2128 60 2162 94
rect 2196 60 2230 94
rect 2264 60 2298 94
rect 2498 60 2532 94
rect 2566 60 2600 94
rect 2634 60 2668 94
rect 2702 60 2736 94
rect 3060 702 3094 736
rect 3128 702 3162 736
rect 3196 702 3230 736
rect 3264 702 3298 736
rect 3498 702 3532 736
rect 3566 702 3600 736
rect 3634 702 3668 736
rect 3702 702 3736 736
rect 3060 634 3094 668
rect 3702 634 3736 668
rect 3060 566 3094 600
rect 3060 498 3094 532
rect 3060 264 3094 298
rect 3060 196 3094 230
rect 3702 566 3736 600
rect 3702 498 3736 532
rect 3702 264 3736 298
rect 3702 196 3736 230
rect 3060 128 3094 162
rect 3702 128 3736 162
rect 3060 60 3094 94
rect 3128 60 3162 94
rect 3196 60 3230 94
rect 3264 60 3298 94
rect 3498 60 3532 94
rect 3566 60 3600 94
rect 3634 60 3668 94
rect 3702 60 3736 94
rect -3940 -298 -3906 -264
rect -3872 -298 -3838 -264
rect -3804 -298 -3770 -264
rect -3736 -298 -3702 -264
rect -3502 -298 -3468 -264
rect -3434 -298 -3400 -264
rect -3366 -298 -3332 -264
rect -3298 -298 -3264 -264
rect -3940 -366 -3906 -332
rect -3298 -366 -3264 -332
rect -3940 -434 -3906 -400
rect -3940 -502 -3906 -468
rect -3940 -736 -3906 -702
rect -3940 -804 -3906 -770
rect -3298 -434 -3264 -400
rect -3298 -502 -3264 -468
rect -3298 -736 -3264 -702
rect -3298 -804 -3264 -770
rect -3940 -872 -3906 -838
rect -3298 -872 -3264 -838
rect -3940 -940 -3906 -906
rect -3872 -940 -3838 -906
rect -3804 -940 -3770 -906
rect -3736 -940 -3702 -906
rect -3502 -940 -3468 -906
rect -3434 -940 -3400 -906
rect -3366 -940 -3332 -906
rect -3298 -940 -3264 -906
rect -2940 -298 -2906 -264
rect -2872 -298 -2838 -264
rect -2804 -298 -2770 -264
rect -2736 -298 -2702 -264
rect -2502 -298 -2468 -264
rect -2434 -298 -2400 -264
rect -2366 -298 -2332 -264
rect -2298 -298 -2264 -264
rect -2940 -366 -2906 -332
rect -2298 -366 -2264 -332
rect -2940 -434 -2906 -400
rect -2940 -502 -2906 -468
rect -2940 -736 -2906 -702
rect -2940 -804 -2906 -770
rect -2298 -434 -2264 -400
rect -2298 -502 -2264 -468
rect -2298 -736 -2264 -702
rect -2298 -804 -2264 -770
rect -2940 -872 -2906 -838
rect -2298 -872 -2264 -838
rect -2940 -940 -2906 -906
rect -2872 -940 -2838 -906
rect -2804 -940 -2770 -906
rect -2736 -940 -2702 -906
rect -2502 -940 -2468 -906
rect -2434 -940 -2400 -906
rect -2366 -940 -2332 -906
rect -2298 -940 -2264 -906
rect -1940 -298 -1906 -264
rect -1872 -298 -1838 -264
rect -1804 -298 -1770 -264
rect -1736 -298 -1702 -264
rect -1502 -298 -1468 -264
rect -1434 -298 -1400 -264
rect -1366 -298 -1332 -264
rect -1298 -298 -1264 -264
rect -1940 -366 -1906 -332
rect -1298 -366 -1264 -332
rect -1940 -434 -1906 -400
rect -1940 -502 -1906 -468
rect -1940 -736 -1906 -702
rect -1940 -804 -1906 -770
rect -1298 -434 -1264 -400
rect -1298 -502 -1264 -468
rect -1298 -736 -1264 -702
rect -1298 -804 -1264 -770
rect -1940 -872 -1906 -838
rect -1298 -872 -1264 -838
rect -1940 -940 -1906 -906
rect -1872 -940 -1838 -906
rect -1804 -940 -1770 -906
rect -1736 -940 -1702 -906
rect -1502 -940 -1468 -906
rect -1434 -940 -1400 -906
rect -1366 -940 -1332 -906
rect -1298 -940 -1264 -906
rect -940 -298 -906 -264
rect -872 -298 -838 -264
rect -804 -298 -770 -264
rect -736 -298 -702 -264
rect -502 -298 -468 -264
rect -434 -298 -400 -264
rect -366 -298 -332 -264
rect -298 -298 -264 -264
rect -940 -366 -906 -332
rect -298 -366 -264 -332
rect -940 -434 -906 -400
rect -940 -502 -906 -468
rect -940 -736 -906 -702
rect -940 -804 -906 -770
rect -298 -434 -264 -400
rect -298 -502 -264 -468
rect -298 -736 -264 -702
rect -298 -804 -264 -770
rect -940 -872 -906 -838
rect -298 -872 -264 -838
rect -940 -940 -906 -906
rect -872 -940 -838 -906
rect -804 -940 -770 -906
rect -736 -940 -702 -906
rect -502 -940 -468 -906
rect -434 -940 -400 -906
rect -366 -940 -332 -906
rect -298 -940 -264 -906
rect 60 -298 94 -264
rect 128 -298 162 -264
rect 196 -298 230 -264
rect 264 -298 298 -264
rect 498 -298 532 -264
rect 566 -298 600 -264
rect 634 -298 668 -264
rect 702 -298 736 -264
rect 60 -366 94 -332
rect 702 -366 736 -332
rect 60 -434 94 -400
rect 60 -502 94 -468
rect 60 -736 94 -702
rect 60 -804 94 -770
rect 702 -434 736 -400
rect 702 -502 736 -468
rect 702 -736 736 -702
rect 702 -804 736 -770
rect 60 -872 94 -838
rect 702 -872 736 -838
rect 60 -940 94 -906
rect 128 -940 162 -906
rect 196 -940 230 -906
rect 264 -940 298 -906
rect 498 -940 532 -906
rect 566 -940 600 -906
rect 634 -940 668 -906
rect 702 -940 736 -906
rect 1060 -298 1094 -264
rect 1128 -298 1162 -264
rect 1196 -298 1230 -264
rect 1264 -298 1298 -264
rect 1498 -298 1532 -264
rect 1566 -298 1600 -264
rect 1634 -298 1668 -264
rect 1702 -298 1736 -264
rect 1060 -366 1094 -332
rect 1702 -366 1736 -332
rect 1060 -434 1094 -400
rect 1060 -502 1094 -468
rect 1060 -736 1094 -702
rect 1060 -804 1094 -770
rect 1702 -434 1736 -400
rect 1702 -502 1736 -468
rect 1702 -736 1736 -702
rect 1702 -804 1736 -770
rect 1060 -872 1094 -838
rect 1702 -872 1736 -838
rect 1060 -940 1094 -906
rect 1128 -940 1162 -906
rect 1196 -940 1230 -906
rect 1264 -940 1298 -906
rect 1498 -940 1532 -906
rect 1566 -940 1600 -906
rect 1634 -940 1668 -906
rect 1702 -940 1736 -906
rect 2060 -298 2094 -264
rect 2128 -298 2162 -264
rect 2196 -298 2230 -264
rect 2264 -298 2298 -264
rect 2498 -298 2532 -264
rect 2566 -298 2600 -264
rect 2634 -298 2668 -264
rect 2702 -298 2736 -264
rect 2060 -366 2094 -332
rect 2702 -366 2736 -332
rect 2060 -434 2094 -400
rect 2060 -502 2094 -468
rect 2060 -736 2094 -702
rect 2060 -804 2094 -770
rect 2702 -434 2736 -400
rect 2702 -502 2736 -468
rect 2702 -736 2736 -702
rect 2702 -804 2736 -770
rect 2060 -872 2094 -838
rect 2702 -872 2736 -838
rect 2060 -940 2094 -906
rect 2128 -940 2162 -906
rect 2196 -940 2230 -906
rect 2264 -940 2298 -906
rect 2498 -940 2532 -906
rect 2566 -940 2600 -906
rect 2634 -940 2668 -906
rect 2702 -940 2736 -906
rect 3060 -298 3094 -264
rect 3128 -298 3162 -264
rect 3196 -298 3230 -264
rect 3264 -298 3298 -264
rect 3498 -298 3532 -264
rect 3566 -298 3600 -264
rect 3634 -298 3668 -264
rect 3702 -298 3736 -264
rect 3060 -366 3094 -332
rect 3702 -366 3736 -332
rect 3060 -434 3094 -400
rect 3060 -502 3094 -468
rect 3060 -736 3094 -702
rect 3060 -804 3094 -770
rect 3702 -434 3736 -400
rect 3702 -502 3736 -468
rect 3702 -736 3736 -702
rect 3702 -804 3736 -770
rect 3060 -872 3094 -838
rect 3702 -872 3736 -838
rect 3060 -940 3094 -906
rect 3128 -940 3162 -906
rect 3196 -940 3230 -906
rect 3264 -940 3298 -906
rect 3498 -940 3532 -906
rect 3566 -940 3600 -906
rect 3634 -940 3668 -906
rect 3702 -940 3736 -906
rect -940 -1298 -906 -1264
rect -872 -1298 -838 -1264
rect -804 -1298 -770 -1264
rect -736 -1298 -702 -1264
rect -502 -1298 -468 -1264
rect -434 -1298 -400 -1264
rect -366 -1298 -332 -1264
rect -298 -1298 -264 -1264
rect -940 -1366 -906 -1332
rect -298 -1366 -264 -1332
rect -940 -1434 -906 -1400
rect -940 -1502 -906 -1468
rect -940 -1736 -906 -1702
rect -940 -1804 -906 -1770
rect -298 -1434 -264 -1400
rect -298 -1502 -264 -1468
rect -298 -1736 -264 -1702
rect -298 -1804 -264 -1770
rect -940 -1872 -906 -1838
rect -298 -1872 -264 -1838
rect -940 -1940 -906 -1906
rect -872 -1940 -838 -1906
rect -804 -1940 -770 -1906
rect -736 -1940 -702 -1906
rect -502 -1940 -468 -1906
rect -434 -1940 -400 -1906
rect -366 -1940 -332 -1906
rect -298 -1940 -264 -1906
rect 60 -1298 94 -1264
rect 128 -1298 162 -1264
rect 196 -1298 230 -1264
rect 264 -1298 298 -1264
rect 498 -1298 532 -1264
rect 566 -1298 600 -1264
rect 634 -1298 668 -1264
rect 702 -1298 736 -1264
rect 60 -1366 94 -1332
rect 702 -1366 736 -1332
rect 60 -1434 94 -1400
rect 60 -1502 94 -1468
rect 60 -1736 94 -1702
rect 60 -1804 94 -1770
rect 702 -1434 736 -1400
rect 702 -1502 736 -1468
rect 702 -1736 736 -1702
rect 702 -1804 736 -1770
rect 60 -1872 94 -1838
rect 702 -1872 736 -1838
rect 60 -1940 94 -1906
rect 128 -1940 162 -1906
rect 196 -1940 230 -1906
rect 264 -1940 298 -1906
rect 498 -1940 532 -1906
rect 566 -1940 600 -1906
rect 634 -1940 668 -1906
rect 702 -1940 736 -1906
rect 1060 -1298 1094 -1264
rect 1128 -1298 1162 -1264
rect 1196 -1298 1230 -1264
rect 1264 -1298 1298 -1264
rect 1498 -1298 1532 -1264
rect 1566 -1298 1600 -1264
rect 1634 -1298 1668 -1264
rect 1702 -1298 1736 -1264
rect 1060 -1366 1094 -1332
rect 1702 -1366 1736 -1332
rect 1060 -1434 1094 -1400
rect 1060 -1502 1094 -1468
rect 1060 -1736 1094 -1702
rect 1060 -1804 1094 -1770
rect 1702 -1434 1736 -1400
rect 1702 -1502 1736 -1468
rect 1702 -1736 1736 -1702
rect 1702 -1804 1736 -1770
rect 1060 -1872 1094 -1838
rect 1702 -1872 1736 -1838
rect 1060 -1940 1094 -1906
rect 1128 -1940 1162 -1906
rect 1196 -1940 1230 -1906
rect 1264 -1940 1298 -1906
rect 1498 -1940 1532 -1906
rect 1566 -1940 1600 -1906
rect 1634 -1940 1668 -1906
rect 1702 -1940 1736 -1906
rect 2060 -1298 2094 -1264
rect 2128 -1298 2162 -1264
rect 2196 -1298 2230 -1264
rect 2264 -1298 2298 -1264
rect 2498 -1298 2532 -1264
rect 2566 -1298 2600 -1264
rect 2634 -1298 2668 -1264
rect 2702 -1298 2736 -1264
rect 2060 -1366 2094 -1332
rect 2702 -1366 2736 -1332
rect 2060 -1434 2094 -1400
rect 2060 -1502 2094 -1468
rect 2060 -1736 2094 -1702
rect 2060 -1804 2094 -1770
rect 2702 -1434 2736 -1400
rect 2702 -1502 2736 -1468
rect 2702 -1736 2736 -1702
rect 2702 -1804 2736 -1770
rect 2060 -1872 2094 -1838
rect 2702 -1872 2736 -1838
rect 2060 -1940 2094 -1906
rect 2128 -1940 2162 -1906
rect 2196 -1940 2230 -1906
rect 2264 -1940 2298 -1906
rect 2498 -1940 2532 -1906
rect 2566 -1940 2600 -1906
rect 2634 -1940 2668 -1906
rect 2702 -1940 2736 -1906
rect 3060 -1298 3094 -1264
rect 3128 -1298 3162 -1264
rect 3196 -1298 3230 -1264
rect 3264 -1298 3298 -1264
rect 3498 -1298 3532 -1264
rect 3566 -1298 3600 -1264
rect 3634 -1298 3668 -1264
rect 3702 -1298 3736 -1264
rect 3060 -1366 3094 -1332
rect 3702 -1366 3736 -1332
rect 3060 -1434 3094 -1400
rect 3060 -1502 3094 -1468
rect 3060 -1736 3094 -1702
rect 3060 -1804 3094 -1770
rect 3702 -1434 3736 -1400
rect 3702 -1502 3736 -1468
rect 3702 -1736 3736 -1702
rect 3702 -1804 3736 -1770
rect 3060 -1872 3094 -1838
rect 3702 -1872 3736 -1838
rect 3060 -1940 3094 -1906
rect 3128 -1940 3162 -1906
rect 3196 -1940 3230 -1906
rect 3264 -1940 3298 -1906
rect 3498 -1940 3532 -1906
rect 3566 -1940 3600 -1906
rect 3634 -1940 3668 -1906
rect 3702 -1940 3736 -1906
rect -940 -2298 -906 -2264
rect -872 -2298 -838 -2264
rect -804 -2298 -770 -2264
rect -736 -2298 -702 -2264
rect -502 -2298 -468 -2264
rect -434 -2298 -400 -2264
rect -366 -2298 -332 -2264
rect -298 -2298 -264 -2264
rect -940 -2366 -906 -2332
rect -298 -2366 -264 -2332
rect -940 -2434 -906 -2400
rect -940 -2502 -906 -2468
rect -940 -2736 -906 -2702
rect -940 -2804 -906 -2770
rect -298 -2434 -264 -2400
rect -298 -2502 -264 -2468
rect -298 -2736 -264 -2702
rect -298 -2804 -264 -2770
rect -940 -2872 -906 -2838
rect -298 -2872 -264 -2838
rect -940 -2940 -906 -2906
rect -872 -2940 -838 -2906
rect -804 -2940 -770 -2906
rect -736 -2940 -702 -2906
rect -502 -2940 -468 -2906
rect -434 -2940 -400 -2906
rect -366 -2940 -332 -2906
rect -298 -2940 -264 -2906
rect 60 -2298 94 -2264
rect 128 -2298 162 -2264
rect 196 -2298 230 -2264
rect 264 -2298 298 -2264
rect 498 -2298 532 -2264
rect 566 -2298 600 -2264
rect 634 -2298 668 -2264
rect 702 -2298 736 -2264
rect 60 -2366 94 -2332
rect 702 -2366 736 -2332
rect 60 -2434 94 -2400
rect 60 -2502 94 -2468
rect 60 -2736 94 -2702
rect 60 -2804 94 -2770
rect 702 -2434 736 -2400
rect 702 -2502 736 -2468
rect 702 -2736 736 -2702
rect 702 -2804 736 -2770
rect 60 -2872 94 -2838
rect 702 -2872 736 -2838
rect 60 -2940 94 -2906
rect 128 -2940 162 -2906
rect 196 -2940 230 -2906
rect 264 -2940 298 -2906
rect 498 -2940 532 -2906
rect 566 -2940 600 -2906
rect 634 -2940 668 -2906
rect 702 -2940 736 -2906
rect 1060 -2298 1094 -2264
rect 1128 -2298 1162 -2264
rect 1196 -2298 1230 -2264
rect 1264 -2298 1298 -2264
rect 1498 -2298 1532 -2264
rect 1566 -2298 1600 -2264
rect 1634 -2298 1668 -2264
rect 1702 -2298 1736 -2264
rect 1060 -2366 1094 -2332
rect 1702 -2366 1736 -2332
rect 1060 -2434 1094 -2400
rect 1060 -2502 1094 -2468
rect 1060 -2736 1094 -2702
rect 1060 -2804 1094 -2770
rect 1702 -2434 1736 -2400
rect 1702 -2502 1736 -2468
rect 1702 -2736 1736 -2702
rect 1702 -2804 1736 -2770
rect 1060 -2872 1094 -2838
rect 1702 -2872 1736 -2838
rect 1060 -2940 1094 -2906
rect 1128 -2940 1162 -2906
rect 1196 -2940 1230 -2906
rect 1264 -2940 1298 -2906
rect 1498 -2940 1532 -2906
rect 1566 -2940 1600 -2906
rect 1634 -2940 1668 -2906
rect 1702 -2940 1736 -2906
rect 2060 -2298 2094 -2264
rect 2128 -2298 2162 -2264
rect 2196 -2298 2230 -2264
rect 2264 -2298 2298 -2264
rect 2498 -2298 2532 -2264
rect 2566 -2298 2600 -2264
rect 2634 -2298 2668 -2264
rect 2702 -2298 2736 -2264
rect 2060 -2366 2094 -2332
rect 2702 -2366 2736 -2332
rect 2060 -2434 2094 -2400
rect 2060 -2502 2094 -2468
rect 2060 -2736 2094 -2702
rect 2060 -2804 2094 -2770
rect 2702 -2434 2736 -2400
rect 2702 -2502 2736 -2468
rect 2702 -2736 2736 -2702
rect 2702 -2804 2736 -2770
rect 2060 -2872 2094 -2838
rect 2702 -2872 2736 -2838
rect 2060 -2940 2094 -2906
rect 2128 -2940 2162 -2906
rect 2196 -2940 2230 -2906
rect 2264 -2940 2298 -2906
rect 2498 -2940 2532 -2906
rect 2566 -2940 2600 -2906
rect 2634 -2940 2668 -2906
rect 2702 -2940 2736 -2906
rect 3060 -2298 3094 -2264
rect 3128 -2298 3162 -2264
rect 3196 -2298 3230 -2264
rect 3264 -2298 3298 -2264
rect 3498 -2298 3532 -2264
rect 3566 -2298 3600 -2264
rect 3634 -2298 3668 -2264
rect 3702 -2298 3736 -2264
rect 3060 -2366 3094 -2332
rect 3702 -2366 3736 -2332
rect 3060 -2434 3094 -2400
rect 3060 -2502 3094 -2468
rect 3060 -2736 3094 -2702
rect 3060 -2804 3094 -2770
rect 3702 -2434 3736 -2400
rect 3702 -2502 3736 -2468
rect 3702 -2736 3736 -2702
rect 3702 -2804 3736 -2770
rect 3060 -2872 3094 -2838
rect 3702 -2872 3736 -2838
rect 3060 -2940 3094 -2906
rect 3128 -2940 3162 -2906
rect 3196 -2940 3230 -2906
rect 3264 -2940 3298 -2906
rect 3498 -2940 3532 -2906
rect 3566 -2940 3600 -2906
rect 3634 -2940 3668 -2906
rect 3702 -2940 3736 -2906
<< nsubdiffcont >>
rect -3787 1549 -3753 1583
rect -3719 1549 -3685 1583
rect -3519 1549 -3485 1583
rect -3451 1549 -3417 1583
rect -3787 1481 -3753 1515
rect -3451 1481 -3417 1515
rect -3787 1281 -3753 1315
rect -3451 1281 -3417 1315
rect -3787 1213 -3753 1247
rect -3719 1213 -3685 1247
rect -3519 1213 -3485 1247
rect -3451 1213 -3417 1247
rect -2787 1549 -2753 1583
rect -2719 1549 -2685 1583
rect -2519 1549 -2485 1583
rect -2451 1549 -2417 1583
rect -2787 1481 -2753 1515
rect -2451 1481 -2417 1515
rect -2787 1281 -2753 1315
rect -2451 1281 -2417 1315
rect -2787 1213 -2753 1247
rect -2719 1213 -2685 1247
rect -2519 1213 -2485 1247
rect -2451 1213 -2417 1247
rect -1787 1549 -1753 1583
rect -1719 1549 -1685 1583
rect -1519 1549 -1485 1583
rect -1451 1549 -1417 1583
rect -1787 1481 -1753 1515
rect -1451 1481 -1417 1515
rect -1787 1281 -1753 1315
rect -1451 1281 -1417 1315
rect -1787 1213 -1753 1247
rect -1719 1213 -1685 1247
rect -1519 1213 -1485 1247
rect -1451 1213 -1417 1247
rect -787 1549 -753 1583
rect -719 1549 -685 1583
rect -519 1549 -485 1583
rect -451 1549 -417 1583
rect -787 1481 -753 1515
rect -451 1481 -417 1515
rect -787 1281 -753 1315
rect -451 1281 -417 1315
rect -787 1213 -753 1247
rect -719 1213 -685 1247
rect -519 1213 -485 1247
rect -451 1213 -417 1247
rect 213 1549 247 1583
rect 281 1549 315 1583
rect 481 1549 515 1583
rect 549 1549 583 1583
rect 213 1481 247 1515
rect 549 1481 583 1515
rect 213 1281 247 1315
rect 549 1281 583 1315
rect 213 1213 247 1247
rect 281 1213 315 1247
rect 481 1213 515 1247
rect 549 1213 583 1247
rect 1213 1549 1247 1583
rect 1281 1549 1315 1583
rect 1481 1549 1515 1583
rect 1549 1549 1583 1583
rect 1213 1481 1247 1515
rect 1549 1481 1583 1515
rect 1213 1281 1247 1315
rect 1549 1281 1583 1315
rect 1213 1213 1247 1247
rect 1281 1213 1315 1247
rect 1481 1213 1515 1247
rect 1549 1213 1583 1247
rect 2213 1549 2247 1583
rect 2281 1549 2315 1583
rect 2481 1549 2515 1583
rect 2549 1549 2583 1583
rect 2213 1481 2247 1515
rect 2549 1481 2583 1515
rect 2213 1281 2247 1315
rect 2549 1281 2583 1315
rect 2213 1213 2247 1247
rect 2281 1213 2315 1247
rect 2481 1213 2515 1247
rect 2549 1213 2583 1247
rect 3213 1549 3247 1583
rect 3281 1549 3315 1583
rect 3481 1549 3515 1583
rect 3549 1549 3583 1583
rect 3213 1481 3247 1515
rect 3549 1481 3583 1515
rect 3213 1281 3247 1315
rect 3549 1281 3583 1315
rect 3213 1213 3247 1247
rect 3281 1213 3315 1247
rect 3481 1213 3515 1247
rect 3549 1213 3583 1247
rect -3787 549 -3753 583
rect -3719 549 -3685 583
rect -3519 549 -3485 583
rect -3451 549 -3417 583
rect -3787 481 -3753 515
rect -3451 481 -3417 515
rect -3787 281 -3753 315
rect -3451 281 -3417 315
rect -3787 213 -3753 247
rect -3719 213 -3685 247
rect -3519 213 -3485 247
rect -3451 213 -3417 247
rect -2787 549 -2753 583
rect -2719 549 -2685 583
rect -2519 549 -2485 583
rect -2451 549 -2417 583
rect -2787 481 -2753 515
rect -2451 481 -2417 515
rect -2787 281 -2753 315
rect -2451 281 -2417 315
rect -2787 213 -2753 247
rect -2719 213 -2685 247
rect -2519 213 -2485 247
rect -2451 213 -2417 247
rect -1787 549 -1753 583
rect -1719 549 -1685 583
rect -1519 549 -1485 583
rect -1451 549 -1417 583
rect -1787 481 -1753 515
rect -1451 481 -1417 515
rect -1787 281 -1753 315
rect -1451 281 -1417 315
rect -1787 213 -1753 247
rect -1719 213 -1685 247
rect -1519 213 -1485 247
rect -1451 213 -1417 247
rect -787 549 -753 583
rect -719 549 -685 583
rect -519 549 -485 583
rect -451 549 -417 583
rect -787 481 -753 515
rect -451 481 -417 515
rect -787 281 -753 315
rect -451 281 -417 315
rect -787 213 -753 247
rect -719 213 -685 247
rect -519 213 -485 247
rect -451 213 -417 247
rect 1213 549 1247 583
rect 1281 549 1315 583
rect 1481 549 1515 583
rect 1549 549 1583 583
rect 1213 481 1247 515
rect 1549 481 1583 515
rect 1213 281 1247 315
rect 1549 281 1583 315
rect 1213 213 1247 247
rect 1281 213 1315 247
rect 1481 213 1515 247
rect 1549 213 1583 247
rect 2213 549 2247 583
rect 2281 549 2315 583
rect 2481 549 2515 583
rect 2549 549 2583 583
rect 2213 481 2247 515
rect 2549 481 2583 515
rect 2213 281 2247 315
rect 2549 281 2583 315
rect 2213 213 2247 247
rect 2281 213 2315 247
rect 2481 213 2515 247
rect 2549 213 2583 247
rect 3213 549 3247 583
rect 3281 549 3315 583
rect 3481 549 3515 583
rect 3549 549 3583 583
rect 3213 481 3247 515
rect 3549 481 3583 515
rect 3213 281 3247 315
rect 3549 281 3583 315
rect 3213 213 3247 247
rect 3281 213 3315 247
rect 3481 213 3515 247
rect 3549 213 3583 247
rect -3787 -451 -3753 -417
rect -3719 -451 -3685 -417
rect -3519 -451 -3485 -417
rect -3451 -451 -3417 -417
rect -3787 -519 -3753 -485
rect -3451 -519 -3417 -485
rect -3787 -719 -3753 -685
rect -3451 -719 -3417 -685
rect -3787 -787 -3753 -753
rect -3719 -787 -3685 -753
rect -3519 -787 -3485 -753
rect -3451 -787 -3417 -753
rect -2787 -451 -2753 -417
rect -2719 -451 -2685 -417
rect -2519 -451 -2485 -417
rect -2451 -451 -2417 -417
rect -2787 -519 -2753 -485
rect -2451 -519 -2417 -485
rect -2787 -719 -2753 -685
rect -2451 -719 -2417 -685
rect -2787 -787 -2753 -753
rect -2719 -787 -2685 -753
rect -2519 -787 -2485 -753
rect -2451 -787 -2417 -753
rect -1787 -451 -1753 -417
rect -1719 -451 -1685 -417
rect -1519 -451 -1485 -417
rect -1451 -451 -1417 -417
rect -1787 -519 -1753 -485
rect -1451 -519 -1417 -485
rect -1787 -719 -1753 -685
rect -1451 -719 -1417 -685
rect -1787 -787 -1753 -753
rect -1719 -787 -1685 -753
rect -1519 -787 -1485 -753
rect -1451 -787 -1417 -753
rect -787 -451 -753 -417
rect -719 -451 -685 -417
rect -519 -451 -485 -417
rect -451 -451 -417 -417
rect -787 -519 -753 -485
rect -451 -519 -417 -485
rect -787 -719 -753 -685
rect -451 -719 -417 -685
rect -787 -787 -753 -753
rect -719 -787 -685 -753
rect -519 -787 -485 -753
rect -451 -787 -417 -753
rect 213 -451 247 -417
rect 281 -451 315 -417
rect 481 -451 515 -417
rect 549 -451 583 -417
rect 213 -519 247 -485
rect 549 -519 583 -485
rect 213 -719 247 -685
rect 549 -719 583 -685
rect 213 -787 247 -753
rect 281 -787 315 -753
rect 481 -787 515 -753
rect 549 -787 583 -753
rect 1213 -451 1247 -417
rect 1281 -451 1315 -417
rect 1481 -451 1515 -417
rect 1549 -451 1583 -417
rect 1213 -519 1247 -485
rect 1549 -519 1583 -485
rect 1213 -719 1247 -685
rect 1549 -719 1583 -685
rect 1213 -787 1247 -753
rect 1281 -787 1315 -753
rect 1481 -787 1515 -753
rect 1549 -787 1583 -753
rect 2213 -451 2247 -417
rect 2281 -451 2315 -417
rect 2481 -451 2515 -417
rect 2549 -451 2583 -417
rect 2213 -519 2247 -485
rect 2549 -519 2583 -485
rect 2213 -719 2247 -685
rect 2549 -719 2583 -685
rect 2213 -787 2247 -753
rect 2281 -787 2315 -753
rect 2481 -787 2515 -753
rect 2549 -787 2583 -753
rect 3213 -451 3247 -417
rect 3281 -451 3315 -417
rect 3481 -451 3515 -417
rect 3549 -451 3583 -417
rect 3213 -519 3247 -485
rect 3549 -519 3583 -485
rect 3213 -719 3247 -685
rect 3549 -719 3583 -685
rect 3213 -787 3247 -753
rect 3281 -787 3315 -753
rect 3481 -787 3515 -753
rect 3549 -787 3583 -753
rect -787 -1451 -753 -1417
rect -719 -1451 -685 -1417
rect -519 -1451 -485 -1417
rect -451 -1451 -417 -1417
rect -787 -1519 -753 -1485
rect -451 -1519 -417 -1485
rect -787 -1719 -753 -1685
rect -451 -1719 -417 -1685
rect -787 -1787 -753 -1753
rect -719 -1787 -685 -1753
rect -519 -1787 -485 -1753
rect -451 -1787 -417 -1753
rect 213 -1451 247 -1417
rect 281 -1451 315 -1417
rect 481 -1451 515 -1417
rect 549 -1451 583 -1417
rect 213 -1519 247 -1485
rect 549 -1519 583 -1485
rect 213 -1719 247 -1685
rect 549 -1719 583 -1685
rect 213 -1787 247 -1753
rect 281 -1787 315 -1753
rect 481 -1787 515 -1753
rect 549 -1787 583 -1753
rect 1213 -1451 1247 -1417
rect 1281 -1451 1315 -1417
rect 1481 -1451 1515 -1417
rect 1549 -1451 1583 -1417
rect 1213 -1519 1247 -1485
rect 1549 -1519 1583 -1485
rect 1213 -1719 1247 -1685
rect 1549 -1719 1583 -1685
rect 1213 -1787 1247 -1753
rect 1281 -1787 1315 -1753
rect 1481 -1787 1515 -1753
rect 1549 -1787 1583 -1753
rect 2213 -1451 2247 -1417
rect 2281 -1451 2315 -1417
rect 2481 -1451 2515 -1417
rect 2549 -1451 2583 -1417
rect 2213 -1519 2247 -1485
rect 2549 -1519 2583 -1485
rect 2213 -1719 2247 -1685
rect 2549 -1719 2583 -1685
rect 2213 -1787 2247 -1753
rect 2281 -1787 2315 -1753
rect 2481 -1787 2515 -1753
rect 2549 -1787 2583 -1753
rect 3213 -1451 3247 -1417
rect 3281 -1451 3315 -1417
rect 3481 -1451 3515 -1417
rect 3549 -1451 3583 -1417
rect 3213 -1519 3247 -1485
rect 3549 -1519 3583 -1485
rect 3213 -1719 3247 -1685
rect 3549 -1719 3583 -1685
rect 3213 -1787 3247 -1753
rect 3281 -1787 3315 -1753
rect 3481 -1787 3515 -1753
rect 3549 -1787 3583 -1753
rect -787 -2451 -753 -2417
rect -719 -2451 -685 -2417
rect -519 -2451 -485 -2417
rect -451 -2451 -417 -2417
rect -787 -2519 -753 -2485
rect -451 -2519 -417 -2485
rect -787 -2719 -753 -2685
rect -451 -2719 -417 -2685
rect -787 -2787 -753 -2753
rect -719 -2787 -685 -2753
rect -519 -2787 -485 -2753
rect -451 -2787 -417 -2753
rect 213 -2451 247 -2417
rect 281 -2451 315 -2417
rect 481 -2451 515 -2417
rect 549 -2451 583 -2417
rect 213 -2519 247 -2485
rect 549 -2519 583 -2485
rect 213 -2719 247 -2685
rect 549 -2719 583 -2685
rect 213 -2787 247 -2753
rect 281 -2787 315 -2753
rect 481 -2787 515 -2753
rect 549 -2787 583 -2753
rect 1213 -2451 1247 -2417
rect 1281 -2451 1315 -2417
rect 1481 -2451 1515 -2417
rect 1549 -2451 1583 -2417
rect 1213 -2519 1247 -2485
rect 1549 -2519 1583 -2485
rect 1213 -2719 1247 -2685
rect 1549 -2719 1583 -2685
rect 1213 -2787 1247 -2753
rect 1281 -2787 1315 -2753
rect 1481 -2787 1515 -2753
rect 1549 -2787 1583 -2753
rect 2213 -2451 2247 -2417
rect 2281 -2451 2315 -2417
rect 2481 -2451 2515 -2417
rect 2549 -2451 2583 -2417
rect 2213 -2519 2247 -2485
rect 2549 -2519 2583 -2485
rect 2213 -2719 2247 -2685
rect 2549 -2719 2583 -2685
rect 2213 -2787 2247 -2753
rect 2281 -2787 2315 -2753
rect 2481 -2787 2515 -2753
rect 2549 -2787 2583 -2753
rect 3213 -2451 3247 -2417
rect 3281 -2451 3315 -2417
rect 3481 -2451 3515 -2417
rect 3549 -2451 3583 -2417
rect 3213 -2519 3247 -2485
rect 3549 -2519 3583 -2485
rect 3213 -2719 3247 -2685
rect 3549 -2719 3583 -2685
rect 3213 -2787 3247 -2753
rect 3281 -2787 3315 -2753
rect 3481 -2787 3515 -2753
rect 3549 -2787 3583 -2753
<< locali >>
rect -3974 1736 -3230 1770
rect -3974 1702 -3940 1736
rect -3906 1702 -3872 1736
rect -3838 1702 -3804 1736
rect -3770 1702 -3736 1736
rect -3702 1702 -3502 1736
rect -3468 1702 -3434 1736
rect -3400 1702 -3366 1736
rect -3332 1702 -3298 1736
rect -3264 1702 -3230 1736
rect -3974 1669 -3230 1702
rect -3974 1668 -3873 1669
rect -3974 1634 -3940 1668
rect -3906 1634 -3873 1668
rect -3974 1600 -3873 1634
rect -3331 1668 -3230 1669
rect -3331 1634 -3298 1668
rect -3264 1634 -3230 1668
rect -3974 1566 -3940 1600
rect -3906 1566 -3873 1600
rect -3974 1532 -3873 1566
rect -3974 1498 -3940 1532
rect -3906 1498 -3873 1532
rect -3974 1298 -3873 1498
rect -3974 1264 -3940 1298
rect -3906 1264 -3873 1298
rect -3974 1230 -3873 1264
rect -3974 1196 -3940 1230
rect -3906 1196 -3873 1230
rect -3974 1162 -3873 1196
rect -3811 1583 -3393 1607
rect -3811 1549 -3787 1583
rect -3753 1549 -3719 1583
rect -3685 1549 -3519 1583
rect -3485 1549 -3451 1583
rect -3417 1549 -3393 1583
rect -3811 1535 -3393 1549
rect -3811 1515 -3739 1535
rect -3811 1481 -3787 1515
rect -3753 1481 -3739 1515
rect -3811 1315 -3739 1481
rect -3465 1515 -3393 1535
rect -3465 1481 -3451 1515
rect -3417 1481 -3393 1515
rect -3681 1463 -3523 1477
rect -3681 1429 -3667 1463
rect -3633 1449 -3571 1463
rect -3537 1429 -3523 1463
rect -3681 1367 -3653 1429
rect -3551 1367 -3523 1429
rect -3681 1333 -3667 1367
rect -3633 1333 -3571 1347
rect -3537 1333 -3523 1367
rect -3681 1319 -3523 1333
rect -3811 1281 -3787 1315
rect -3753 1281 -3739 1315
rect -3811 1261 -3739 1281
rect -3465 1315 -3393 1481
rect -3465 1281 -3451 1315
rect -3417 1281 -3393 1315
rect -3465 1261 -3393 1281
rect -3811 1247 -3393 1261
rect -3811 1213 -3787 1247
rect -3753 1213 -3719 1247
rect -3685 1213 -3519 1247
rect -3485 1213 -3451 1247
rect -3417 1213 -3393 1247
rect -3811 1189 -3393 1213
rect -3331 1600 -3230 1634
rect -3331 1566 -3298 1600
rect -3264 1566 -3230 1600
rect -3331 1532 -3230 1566
rect -3331 1498 -3298 1532
rect -3264 1498 -3230 1532
rect -3331 1298 -3230 1498
rect -3331 1264 -3298 1298
rect -3264 1264 -3230 1298
rect -3331 1230 -3230 1264
rect -3331 1196 -3298 1230
rect -3264 1196 -3230 1230
rect -3974 1128 -3940 1162
rect -3906 1128 -3873 1162
rect -3974 1127 -3873 1128
rect -3331 1162 -3230 1196
rect -3331 1128 -3298 1162
rect -3264 1128 -3230 1162
rect -3331 1127 -3230 1128
rect -3974 1094 -3230 1127
rect -3974 1060 -3940 1094
rect -3906 1060 -3872 1094
rect -3838 1060 -3804 1094
rect -3770 1060 -3736 1094
rect -3702 1060 -3502 1094
rect -3468 1060 -3434 1094
rect -3400 1060 -3366 1094
rect -3332 1060 -3298 1094
rect -3264 1060 -3230 1094
rect -3974 1026 -3230 1060
rect -2974 1736 -2230 1770
rect -2974 1702 -2940 1736
rect -2906 1702 -2872 1736
rect -2838 1702 -2804 1736
rect -2770 1702 -2736 1736
rect -2702 1702 -2502 1736
rect -2468 1702 -2434 1736
rect -2400 1702 -2366 1736
rect -2332 1702 -2298 1736
rect -2264 1702 -2230 1736
rect -2974 1669 -2230 1702
rect -2974 1668 -2873 1669
rect -2974 1634 -2940 1668
rect -2906 1634 -2873 1668
rect -2974 1600 -2873 1634
rect -2331 1668 -2230 1669
rect -2331 1634 -2298 1668
rect -2264 1634 -2230 1668
rect -2974 1566 -2940 1600
rect -2906 1566 -2873 1600
rect -2974 1532 -2873 1566
rect -2974 1498 -2940 1532
rect -2906 1498 -2873 1532
rect -2974 1298 -2873 1498
rect -2974 1264 -2940 1298
rect -2906 1264 -2873 1298
rect -2974 1230 -2873 1264
rect -2974 1196 -2940 1230
rect -2906 1196 -2873 1230
rect -2974 1162 -2873 1196
rect -2811 1583 -2393 1607
rect -2811 1549 -2787 1583
rect -2753 1549 -2719 1583
rect -2685 1549 -2519 1583
rect -2485 1549 -2451 1583
rect -2417 1549 -2393 1583
rect -2811 1535 -2393 1549
rect -2811 1515 -2739 1535
rect -2811 1481 -2787 1515
rect -2753 1481 -2739 1515
rect -2811 1315 -2739 1481
rect -2465 1515 -2393 1535
rect -2465 1481 -2451 1515
rect -2417 1481 -2393 1515
rect -2681 1463 -2523 1477
rect -2681 1429 -2667 1463
rect -2633 1449 -2571 1463
rect -2537 1429 -2523 1463
rect -2681 1367 -2653 1429
rect -2551 1367 -2523 1429
rect -2681 1333 -2667 1367
rect -2633 1333 -2571 1347
rect -2537 1333 -2523 1367
rect -2681 1319 -2523 1333
rect -2811 1281 -2787 1315
rect -2753 1281 -2739 1315
rect -2811 1261 -2739 1281
rect -2465 1315 -2393 1481
rect -2465 1281 -2451 1315
rect -2417 1281 -2393 1315
rect -2465 1261 -2393 1281
rect -2811 1247 -2393 1261
rect -2811 1213 -2787 1247
rect -2753 1213 -2719 1247
rect -2685 1213 -2519 1247
rect -2485 1213 -2451 1247
rect -2417 1213 -2393 1247
rect -2811 1189 -2393 1213
rect -2331 1600 -2230 1634
rect -2331 1566 -2298 1600
rect -2264 1566 -2230 1600
rect -2331 1532 -2230 1566
rect -2331 1498 -2298 1532
rect -2264 1498 -2230 1532
rect -2331 1298 -2230 1498
rect -2331 1264 -2298 1298
rect -2264 1264 -2230 1298
rect -2331 1230 -2230 1264
rect -2331 1196 -2298 1230
rect -2264 1196 -2230 1230
rect -2974 1128 -2940 1162
rect -2906 1128 -2873 1162
rect -2974 1127 -2873 1128
rect -2331 1162 -2230 1196
rect -2331 1128 -2298 1162
rect -2264 1128 -2230 1162
rect -2331 1127 -2230 1128
rect -2974 1094 -2230 1127
rect -2974 1060 -2940 1094
rect -2906 1060 -2872 1094
rect -2838 1060 -2804 1094
rect -2770 1060 -2736 1094
rect -2702 1060 -2502 1094
rect -2468 1060 -2434 1094
rect -2400 1060 -2366 1094
rect -2332 1060 -2298 1094
rect -2264 1060 -2230 1094
rect -2974 1026 -2230 1060
rect -1974 1736 -1230 1770
rect -1974 1702 -1940 1736
rect -1906 1702 -1872 1736
rect -1838 1702 -1804 1736
rect -1770 1702 -1736 1736
rect -1702 1702 -1502 1736
rect -1468 1702 -1434 1736
rect -1400 1702 -1366 1736
rect -1332 1702 -1298 1736
rect -1264 1702 -1230 1736
rect -1974 1669 -1230 1702
rect -1974 1668 -1873 1669
rect -1974 1634 -1940 1668
rect -1906 1634 -1873 1668
rect -1974 1600 -1873 1634
rect -1331 1668 -1230 1669
rect -1331 1634 -1298 1668
rect -1264 1634 -1230 1668
rect -1974 1566 -1940 1600
rect -1906 1566 -1873 1600
rect -1974 1532 -1873 1566
rect -1974 1498 -1940 1532
rect -1906 1498 -1873 1532
rect -1974 1298 -1873 1498
rect -1974 1264 -1940 1298
rect -1906 1264 -1873 1298
rect -1974 1230 -1873 1264
rect -1974 1196 -1940 1230
rect -1906 1196 -1873 1230
rect -1974 1162 -1873 1196
rect -1811 1583 -1393 1607
rect -1811 1549 -1787 1583
rect -1753 1549 -1719 1583
rect -1685 1549 -1519 1583
rect -1485 1549 -1451 1583
rect -1417 1549 -1393 1583
rect -1811 1535 -1393 1549
rect -1811 1515 -1739 1535
rect -1811 1481 -1787 1515
rect -1753 1481 -1739 1515
rect -1811 1315 -1739 1481
rect -1465 1515 -1393 1535
rect -1465 1481 -1451 1515
rect -1417 1481 -1393 1515
rect -1681 1463 -1523 1477
rect -1681 1429 -1667 1463
rect -1633 1449 -1571 1463
rect -1537 1429 -1523 1463
rect -1681 1367 -1653 1429
rect -1551 1367 -1523 1429
rect -1681 1333 -1667 1367
rect -1633 1333 -1571 1347
rect -1537 1333 -1523 1367
rect -1681 1319 -1523 1333
rect -1811 1281 -1787 1315
rect -1753 1281 -1739 1315
rect -1811 1261 -1739 1281
rect -1465 1315 -1393 1481
rect -1465 1281 -1451 1315
rect -1417 1281 -1393 1315
rect -1465 1261 -1393 1281
rect -1811 1247 -1393 1261
rect -1811 1213 -1787 1247
rect -1753 1213 -1719 1247
rect -1685 1213 -1519 1247
rect -1485 1213 -1451 1247
rect -1417 1213 -1393 1247
rect -1811 1189 -1393 1213
rect -1331 1600 -1230 1634
rect -1331 1566 -1298 1600
rect -1264 1566 -1230 1600
rect -1331 1532 -1230 1566
rect -1331 1498 -1298 1532
rect -1264 1498 -1230 1532
rect -1331 1298 -1230 1498
rect -1331 1264 -1298 1298
rect -1264 1264 -1230 1298
rect -1331 1230 -1230 1264
rect -1331 1196 -1298 1230
rect -1264 1196 -1230 1230
rect -1974 1128 -1940 1162
rect -1906 1128 -1873 1162
rect -1974 1127 -1873 1128
rect -1331 1162 -1230 1196
rect -1331 1128 -1298 1162
rect -1264 1128 -1230 1162
rect -1331 1127 -1230 1128
rect -1974 1094 -1230 1127
rect -1974 1060 -1940 1094
rect -1906 1060 -1872 1094
rect -1838 1060 -1804 1094
rect -1770 1060 -1736 1094
rect -1702 1060 -1502 1094
rect -1468 1060 -1434 1094
rect -1400 1060 -1366 1094
rect -1332 1060 -1298 1094
rect -1264 1060 -1230 1094
rect -1974 1026 -1230 1060
rect -974 1736 -230 1770
rect -974 1702 -940 1736
rect -906 1702 -872 1736
rect -838 1702 -804 1736
rect -770 1702 -736 1736
rect -702 1702 -502 1736
rect -468 1702 -434 1736
rect -400 1702 -366 1736
rect -332 1702 -298 1736
rect -264 1702 -230 1736
rect -974 1669 -230 1702
rect -974 1668 -873 1669
rect -974 1634 -940 1668
rect -906 1634 -873 1668
rect -974 1600 -873 1634
rect -331 1668 -230 1669
rect -331 1634 -298 1668
rect -264 1634 -230 1668
rect -974 1566 -940 1600
rect -906 1566 -873 1600
rect -974 1532 -873 1566
rect -974 1498 -940 1532
rect -906 1498 -873 1532
rect -974 1298 -873 1498
rect -974 1264 -940 1298
rect -906 1264 -873 1298
rect -974 1230 -873 1264
rect -974 1196 -940 1230
rect -906 1196 -873 1230
rect -974 1162 -873 1196
rect -811 1583 -393 1607
rect -811 1549 -787 1583
rect -753 1549 -719 1583
rect -685 1549 -519 1583
rect -485 1549 -451 1583
rect -417 1549 -393 1583
rect -811 1535 -393 1549
rect -811 1515 -739 1535
rect -811 1481 -787 1515
rect -753 1481 -739 1515
rect -811 1315 -739 1481
rect -465 1515 -393 1535
rect -465 1481 -451 1515
rect -417 1481 -393 1515
rect -681 1463 -523 1477
rect -681 1429 -667 1463
rect -633 1449 -571 1463
rect -537 1429 -523 1463
rect -681 1367 -653 1429
rect -551 1367 -523 1429
rect -681 1333 -667 1367
rect -633 1333 -571 1347
rect -537 1333 -523 1367
rect -681 1319 -523 1333
rect -811 1281 -787 1315
rect -753 1281 -739 1315
rect -811 1261 -739 1281
rect -465 1315 -393 1481
rect -465 1281 -451 1315
rect -417 1281 -393 1315
rect -465 1261 -393 1281
rect -811 1247 -393 1261
rect -811 1213 -787 1247
rect -753 1213 -719 1247
rect -685 1213 -519 1247
rect -485 1213 -451 1247
rect -417 1213 -393 1247
rect -811 1189 -393 1213
rect -331 1600 -230 1634
rect -331 1566 -298 1600
rect -264 1566 -230 1600
rect -331 1532 -230 1566
rect -331 1498 -298 1532
rect -264 1498 -230 1532
rect -331 1298 -230 1498
rect -331 1264 -298 1298
rect -264 1264 -230 1298
rect -331 1230 -230 1264
rect -331 1196 -298 1230
rect -264 1196 -230 1230
rect -974 1128 -940 1162
rect -906 1128 -873 1162
rect -974 1127 -873 1128
rect -331 1162 -230 1196
rect -331 1128 -298 1162
rect -264 1128 -230 1162
rect -331 1127 -230 1128
rect -974 1094 -230 1127
rect -974 1060 -940 1094
rect -906 1060 -872 1094
rect -838 1060 -804 1094
rect -770 1060 -736 1094
rect -702 1060 -502 1094
rect -468 1060 -434 1094
rect -400 1060 -366 1094
rect -332 1060 -298 1094
rect -264 1060 -230 1094
rect -974 1026 -230 1060
rect 26 1736 770 1770
rect 26 1702 60 1736
rect 94 1702 128 1736
rect 162 1702 196 1736
rect 230 1702 264 1736
rect 298 1702 498 1736
rect 532 1702 566 1736
rect 600 1702 634 1736
rect 668 1702 702 1736
rect 736 1702 770 1736
rect 26 1669 770 1702
rect 26 1668 127 1669
rect 26 1634 60 1668
rect 94 1634 127 1668
rect 26 1600 127 1634
rect 669 1668 770 1669
rect 669 1634 702 1668
rect 736 1634 770 1668
rect 26 1566 60 1600
rect 94 1566 127 1600
rect 26 1532 127 1566
rect 26 1498 60 1532
rect 94 1498 127 1532
rect 26 1298 127 1498
rect 26 1264 60 1298
rect 94 1264 127 1298
rect 26 1230 127 1264
rect 26 1196 60 1230
rect 94 1196 127 1230
rect 26 1162 127 1196
rect 189 1583 607 1607
rect 189 1549 213 1583
rect 247 1549 281 1583
rect 315 1549 481 1583
rect 515 1549 549 1583
rect 583 1549 607 1583
rect 189 1535 607 1549
rect 189 1515 261 1535
rect 189 1481 213 1515
rect 247 1481 261 1515
rect 189 1315 261 1481
rect 535 1515 607 1535
rect 535 1481 549 1515
rect 583 1481 607 1515
rect 319 1463 477 1477
rect 319 1429 333 1463
rect 367 1449 429 1463
rect 463 1429 477 1463
rect 319 1367 347 1429
rect 449 1367 477 1429
rect 319 1333 333 1367
rect 367 1333 429 1347
rect 463 1333 477 1367
rect 319 1319 477 1333
rect 189 1281 213 1315
rect 247 1281 261 1315
rect 189 1261 261 1281
rect 535 1315 607 1481
rect 535 1281 549 1315
rect 583 1281 607 1315
rect 535 1261 607 1281
rect 189 1247 607 1261
rect 189 1213 213 1247
rect 247 1213 281 1247
rect 315 1213 481 1247
rect 515 1213 549 1247
rect 583 1213 607 1247
rect 189 1189 607 1213
rect 669 1600 770 1634
rect 669 1566 702 1600
rect 736 1566 770 1600
rect 669 1532 770 1566
rect 669 1498 702 1532
rect 736 1498 770 1532
rect 669 1298 770 1498
rect 669 1264 702 1298
rect 736 1264 770 1298
rect 669 1230 770 1264
rect 669 1196 702 1230
rect 736 1196 770 1230
rect 26 1128 60 1162
rect 94 1128 127 1162
rect 26 1127 127 1128
rect 669 1162 770 1196
rect 669 1128 702 1162
rect 736 1128 770 1162
rect 669 1127 770 1128
rect 26 1094 770 1127
rect 26 1060 60 1094
rect 94 1060 128 1094
rect 162 1060 196 1094
rect 230 1060 264 1094
rect 298 1060 498 1094
rect 532 1060 566 1094
rect 600 1060 634 1094
rect 668 1060 702 1094
rect 736 1060 770 1094
rect 26 1026 770 1060
rect 1026 1736 1770 1770
rect 1026 1702 1060 1736
rect 1094 1702 1128 1736
rect 1162 1702 1196 1736
rect 1230 1702 1264 1736
rect 1298 1702 1498 1736
rect 1532 1702 1566 1736
rect 1600 1702 1634 1736
rect 1668 1702 1702 1736
rect 1736 1702 1770 1736
rect 1026 1669 1770 1702
rect 1026 1668 1127 1669
rect 1026 1634 1060 1668
rect 1094 1634 1127 1668
rect 1026 1600 1127 1634
rect 1669 1668 1770 1669
rect 1669 1634 1702 1668
rect 1736 1634 1770 1668
rect 1026 1566 1060 1600
rect 1094 1566 1127 1600
rect 1026 1532 1127 1566
rect 1026 1498 1060 1532
rect 1094 1498 1127 1532
rect 1026 1298 1127 1498
rect 1026 1264 1060 1298
rect 1094 1264 1127 1298
rect 1026 1230 1127 1264
rect 1026 1196 1060 1230
rect 1094 1196 1127 1230
rect 1026 1162 1127 1196
rect 1189 1583 1607 1607
rect 1189 1549 1213 1583
rect 1247 1549 1281 1583
rect 1315 1549 1481 1583
rect 1515 1549 1549 1583
rect 1583 1549 1607 1583
rect 1189 1535 1607 1549
rect 1189 1515 1261 1535
rect 1189 1481 1213 1515
rect 1247 1481 1261 1515
rect 1189 1315 1261 1481
rect 1535 1515 1607 1535
rect 1535 1481 1549 1515
rect 1583 1481 1607 1515
rect 1319 1463 1477 1477
rect 1319 1429 1333 1463
rect 1367 1449 1429 1463
rect 1463 1429 1477 1463
rect 1319 1367 1347 1429
rect 1449 1367 1477 1429
rect 1319 1333 1333 1367
rect 1367 1333 1429 1347
rect 1463 1333 1477 1367
rect 1319 1319 1477 1333
rect 1189 1281 1213 1315
rect 1247 1281 1261 1315
rect 1189 1261 1261 1281
rect 1535 1315 1607 1481
rect 1535 1281 1549 1315
rect 1583 1281 1607 1315
rect 1535 1261 1607 1281
rect 1189 1247 1607 1261
rect 1189 1213 1213 1247
rect 1247 1213 1281 1247
rect 1315 1213 1481 1247
rect 1515 1213 1549 1247
rect 1583 1213 1607 1247
rect 1189 1189 1607 1213
rect 1669 1600 1770 1634
rect 1669 1566 1702 1600
rect 1736 1566 1770 1600
rect 1669 1532 1770 1566
rect 1669 1498 1702 1532
rect 1736 1498 1770 1532
rect 1669 1298 1770 1498
rect 1669 1264 1702 1298
rect 1736 1264 1770 1298
rect 1669 1230 1770 1264
rect 1669 1196 1702 1230
rect 1736 1196 1770 1230
rect 1026 1128 1060 1162
rect 1094 1128 1127 1162
rect 1026 1127 1127 1128
rect 1669 1162 1770 1196
rect 1669 1128 1702 1162
rect 1736 1128 1770 1162
rect 1669 1127 1770 1128
rect 1026 1094 1770 1127
rect 1026 1060 1060 1094
rect 1094 1060 1128 1094
rect 1162 1060 1196 1094
rect 1230 1060 1264 1094
rect 1298 1060 1498 1094
rect 1532 1060 1566 1094
rect 1600 1060 1634 1094
rect 1668 1060 1702 1094
rect 1736 1060 1770 1094
rect 1026 1026 1770 1060
rect 2026 1736 2770 1770
rect 2026 1702 2060 1736
rect 2094 1702 2128 1736
rect 2162 1702 2196 1736
rect 2230 1702 2264 1736
rect 2298 1702 2498 1736
rect 2532 1702 2566 1736
rect 2600 1702 2634 1736
rect 2668 1702 2702 1736
rect 2736 1702 2770 1736
rect 2026 1669 2770 1702
rect 2026 1668 2127 1669
rect 2026 1634 2060 1668
rect 2094 1634 2127 1668
rect 2026 1600 2127 1634
rect 2669 1668 2770 1669
rect 2669 1634 2702 1668
rect 2736 1634 2770 1668
rect 2026 1566 2060 1600
rect 2094 1566 2127 1600
rect 2026 1532 2127 1566
rect 2026 1498 2060 1532
rect 2094 1498 2127 1532
rect 2026 1298 2127 1498
rect 2026 1264 2060 1298
rect 2094 1264 2127 1298
rect 2026 1230 2127 1264
rect 2026 1196 2060 1230
rect 2094 1196 2127 1230
rect 2026 1162 2127 1196
rect 2189 1583 2607 1607
rect 2189 1549 2213 1583
rect 2247 1549 2281 1583
rect 2315 1549 2481 1583
rect 2515 1549 2549 1583
rect 2583 1549 2607 1583
rect 2189 1535 2607 1549
rect 2189 1515 2261 1535
rect 2189 1481 2213 1515
rect 2247 1481 2261 1515
rect 2189 1315 2261 1481
rect 2535 1515 2607 1535
rect 2535 1481 2549 1515
rect 2583 1481 2607 1515
rect 2319 1463 2477 1477
rect 2319 1429 2333 1463
rect 2367 1449 2429 1463
rect 2463 1429 2477 1463
rect 2319 1367 2347 1429
rect 2449 1367 2477 1429
rect 2319 1333 2333 1367
rect 2367 1333 2429 1347
rect 2463 1333 2477 1367
rect 2319 1319 2477 1333
rect 2189 1281 2213 1315
rect 2247 1281 2261 1315
rect 2189 1261 2261 1281
rect 2535 1315 2607 1481
rect 2535 1281 2549 1315
rect 2583 1281 2607 1315
rect 2535 1261 2607 1281
rect 2189 1247 2607 1261
rect 2189 1213 2213 1247
rect 2247 1213 2281 1247
rect 2315 1213 2481 1247
rect 2515 1213 2549 1247
rect 2583 1213 2607 1247
rect 2189 1189 2607 1213
rect 2669 1600 2770 1634
rect 2669 1566 2702 1600
rect 2736 1566 2770 1600
rect 2669 1532 2770 1566
rect 2669 1498 2702 1532
rect 2736 1498 2770 1532
rect 2669 1298 2770 1498
rect 2669 1264 2702 1298
rect 2736 1264 2770 1298
rect 2669 1230 2770 1264
rect 2669 1196 2702 1230
rect 2736 1196 2770 1230
rect 2026 1128 2060 1162
rect 2094 1128 2127 1162
rect 2026 1127 2127 1128
rect 2669 1162 2770 1196
rect 2669 1128 2702 1162
rect 2736 1128 2770 1162
rect 2669 1127 2770 1128
rect 2026 1094 2770 1127
rect 2026 1060 2060 1094
rect 2094 1060 2128 1094
rect 2162 1060 2196 1094
rect 2230 1060 2264 1094
rect 2298 1060 2498 1094
rect 2532 1060 2566 1094
rect 2600 1060 2634 1094
rect 2668 1060 2702 1094
rect 2736 1060 2770 1094
rect 2026 1026 2770 1060
rect 3026 1736 3770 1770
rect 3026 1702 3060 1736
rect 3094 1702 3128 1736
rect 3162 1702 3196 1736
rect 3230 1702 3264 1736
rect 3298 1702 3498 1736
rect 3532 1702 3566 1736
rect 3600 1702 3634 1736
rect 3668 1702 3702 1736
rect 3736 1702 3770 1736
rect 3026 1669 3770 1702
rect 3026 1668 3127 1669
rect 3026 1634 3060 1668
rect 3094 1634 3127 1668
rect 3026 1600 3127 1634
rect 3669 1668 3770 1669
rect 3669 1634 3702 1668
rect 3736 1634 3770 1668
rect 3026 1566 3060 1600
rect 3094 1566 3127 1600
rect 3026 1532 3127 1566
rect 3026 1498 3060 1532
rect 3094 1498 3127 1532
rect 3026 1298 3127 1498
rect 3026 1264 3060 1298
rect 3094 1264 3127 1298
rect 3026 1230 3127 1264
rect 3026 1196 3060 1230
rect 3094 1196 3127 1230
rect 3026 1162 3127 1196
rect 3189 1583 3607 1607
rect 3189 1549 3213 1583
rect 3247 1549 3281 1583
rect 3315 1549 3481 1583
rect 3515 1549 3549 1583
rect 3583 1549 3607 1583
rect 3189 1535 3607 1549
rect 3189 1515 3261 1535
rect 3189 1481 3213 1515
rect 3247 1481 3261 1515
rect 3189 1315 3261 1481
rect 3535 1515 3607 1535
rect 3535 1481 3549 1515
rect 3583 1481 3607 1515
rect 3319 1463 3477 1477
rect 3319 1429 3333 1463
rect 3367 1449 3429 1463
rect 3463 1429 3477 1463
rect 3319 1367 3347 1429
rect 3449 1367 3477 1429
rect 3319 1333 3333 1367
rect 3367 1333 3429 1347
rect 3463 1333 3477 1367
rect 3319 1319 3477 1333
rect 3189 1281 3213 1315
rect 3247 1281 3261 1315
rect 3189 1261 3261 1281
rect 3535 1315 3607 1481
rect 3535 1281 3549 1315
rect 3583 1281 3607 1315
rect 3535 1261 3607 1281
rect 3189 1247 3607 1261
rect 3189 1213 3213 1247
rect 3247 1213 3281 1247
rect 3315 1213 3481 1247
rect 3515 1213 3549 1247
rect 3583 1213 3607 1247
rect 3189 1189 3607 1213
rect 3669 1600 3770 1634
rect 3669 1566 3702 1600
rect 3736 1566 3770 1600
rect 3669 1532 3770 1566
rect 3669 1498 3702 1532
rect 3736 1498 3770 1532
rect 3669 1298 3770 1498
rect 3669 1264 3702 1298
rect 3736 1264 3770 1298
rect 3669 1230 3770 1264
rect 3669 1196 3702 1230
rect 3736 1196 3770 1230
rect 3026 1128 3060 1162
rect 3094 1128 3127 1162
rect 3026 1127 3127 1128
rect 3669 1162 3770 1196
rect 3669 1128 3702 1162
rect 3736 1128 3770 1162
rect 3669 1127 3770 1128
rect 3026 1094 3770 1127
rect 3026 1060 3060 1094
rect 3094 1060 3128 1094
rect 3162 1060 3196 1094
rect 3230 1060 3264 1094
rect 3298 1060 3498 1094
rect 3532 1060 3566 1094
rect 3600 1060 3634 1094
rect 3668 1060 3702 1094
rect 3736 1060 3770 1094
rect 3026 1026 3770 1060
rect -3974 736 -3230 770
rect -3974 702 -3940 736
rect -3906 702 -3872 736
rect -3838 702 -3804 736
rect -3770 702 -3736 736
rect -3702 702 -3502 736
rect -3468 702 -3434 736
rect -3400 702 -3366 736
rect -3332 702 -3298 736
rect -3264 702 -3230 736
rect -3974 669 -3230 702
rect -3974 668 -3873 669
rect -3974 634 -3940 668
rect -3906 634 -3873 668
rect -3974 600 -3873 634
rect -3331 668 -3230 669
rect -3331 634 -3298 668
rect -3264 634 -3230 668
rect -3974 566 -3940 600
rect -3906 566 -3873 600
rect -3974 532 -3873 566
rect -3974 498 -3940 532
rect -3906 498 -3873 532
rect -3974 298 -3873 498
rect -3974 264 -3940 298
rect -3906 264 -3873 298
rect -3974 230 -3873 264
rect -3974 196 -3940 230
rect -3906 196 -3873 230
rect -3974 162 -3873 196
rect -3811 583 -3393 607
rect -3811 549 -3787 583
rect -3753 549 -3719 583
rect -3685 549 -3519 583
rect -3485 549 -3451 583
rect -3417 549 -3393 583
rect -3811 535 -3393 549
rect -3811 515 -3739 535
rect -3811 481 -3787 515
rect -3753 481 -3739 515
rect -3811 315 -3739 481
rect -3465 515 -3393 535
rect -3465 481 -3451 515
rect -3417 481 -3393 515
rect -3681 463 -3523 477
rect -3681 429 -3667 463
rect -3633 449 -3571 463
rect -3537 429 -3523 463
rect -3681 367 -3653 429
rect -3551 367 -3523 429
rect -3681 333 -3667 367
rect -3633 333 -3571 347
rect -3537 333 -3523 367
rect -3681 319 -3523 333
rect -3811 281 -3787 315
rect -3753 281 -3739 315
rect -3811 261 -3739 281
rect -3465 315 -3393 481
rect -3465 281 -3451 315
rect -3417 281 -3393 315
rect -3465 261 -3393 281
rect -3811 247 -3393 261
rect -3811 213 -3787 247
rect -3753 213 -3719 247
rect -3685 213 -3519 247
rect -3485 213 -3451 247
rect -3417 213 -3393 247
rect -3811 189 -3393 213
rect -3331 600 -3230 634
rect -3331 566 -3298 600
rect -3264 566 -3230 600
rect -3331 532 -3230 566
rect -3331 498 -3298 532
rect -3264 498 -3230 532
rect -3331 298 -3230 498
rect -3331 264 -3298 298
rect -3264 264 -3230 298
rect -3331 230 -3230 264
rect -3331 196 -3298 230
rect -3264 196 -3230 230
rect -3974 128 -3940 162
rect -3906 128 -3873 162
rect -3974 127 -3873 128
rect -3331 162 -3230 196
rect -3331 128 -3298 162
rect -3264 128 -3230 162
rect -3331 127 -3230 128
rect -3974 94 -3230 127
rect -3974 60 -3940 94
rect -3906 60 -3872 94
rect -3838 60 -3804 94
rect -3770 60 -3736 94
rect -3702 60 -3502 94
rect -3468 60 -3434 94
rect -3400 60 -3366 94
rect -3332 60 -3298 94
rect -3264 60 -3230 94
rect -3974 26 -3230 60
rect -2974 736 -2230 770
rect -2974 702 -2940 736
rect -2906 702 -2872 736
rect -2838 702 -2804 736
rect -2770 702 -2736 736
rect -2702 702 -2502 736
rect -2468 702 -2434 736
rect -2400 702 -2366 736
rect -2332 702 -2298 736
rect -2264 702 -2230 736
rect -2974 669 -2230 702
rect -2974 668 -2873 669
rect -2974 634 -2940 668
rect -2906 634 -2873 668
rect -2974 600 -2873 634
rect -2331 668 -2230 669
rect -2331 634 -2298 668
rect -2264 634 -2230 668
rect -2974 566 -2940 600
rect -2906 566 -2873 600
rect -2974 532 -2873 566
rect -2974 498 -2940 532
rect -2906 498 -2873 532
rect -2974 298 -2873 498
rect -2974 264 -2940 298
rect -2906 264 -2873 298
rect -2974 230 -2873 264
rect -2974 196 -2940 230
rect -2906 196 -2873 230
rect -2974 162 -2873 196
rect -2811 583 -2393 607
rect -2811 549 -2787 583
rect -2753 549 -2719 583
rect -2685 549 -2519 583
rect -2485 549 -2451 583
rect -2417 549 -2393 583
rect -2811 535 -2393 549
rect -2811 515 -2739 535
rect -2811 481 -2787 515
rect -2753 481 -2739 515
rect -2811 315 -2739 481
rect -2465 515 -2393 535
rect -2465 481 -2451 515
rect -2417 481 -2393 515
rect -2681 463 -2523 477
rect -2681 429 -2667 463
rect -2633 449 -2571 463
rect -2537 429 -2523 463
rect -2681 367 -2653 429
rect -2551 367 -2523 429
rect -2681 333 -2667 367
rect -2633 333 -2571 347
rect -2537 333 -2523 367
rect -2681 319 -2523 333
rect -2811 281 -2787 315
rect -2753 281 -2739 315
rect -2811 261 -2739 281
rect -2465 315 -2393 481
rect -2465 281 -2451 315
rect -2417 281 -2393 315
rect -2465 261 -2393 281
rect -2811 247 -2393 261
rect -2811 213 -2787 247
rect -2753 213 -2719 247
rect -2685 213 -2519 247
rect -2485 213 -2451 247
rect -2417 213 -2393 247
rect -2811 189 -2393 213
rect -2331 600 -2230 634
rect -2331 566 -2298 600
rect -2264 566 -2230 600
rect -2331 532 -2230 566
rect -2331 498 -2298 532
rect -2264 498 -2230 532
rect -2331 298 -2230 498
rect -2331 264 -2298 298
rect -2264 264 -2230 298
rect -2331 230 -2230 264
rect -2331 196 -2298 230
rect -2264 196 -2230 230
rect -2974 128 -2940 162
rect -2906 128 -2873 162
rect -2974 127 -2873 128
rect -2331 162 -2230 196
rect -2331 128 -2298 162
rect -2264 128 -2230 162
rect -2331 127 -2230 128
rect -2974 94 -2230 127
rect -2974 60 -2940 94
rect -2906 60 -2872 94
rect -2838 60 -2804 94
rect -2770 60 -2736 94
rect -2702 60 -2502 94
rect -2468 60 -2434 94
rect -2400 60 -2366 94
rect -2332 60 -2298 94
rect -2264 60 -2230 94
rect -2974 26 -2230 60
rect -1974 736 -1230 770
rect -1974 702 -1940 736
rect -1906 702 -1872 736
rect -1838 702 -1804 736
rect -1770 702 -1736 736
rect -1702 702 -1502 736
rect -1468 702 -1434 736
rect -1400 702 -1366 736
rect -1332 702 -1298 736
rect -1264 702 -1230 736
rect -1974 669 -1230 702
rect -1974 668 -1873 669
rect -1974 634 -1940 668
rect -1906 634 -1873 668
rect -1974 600 -1873 634
rect -1331 668 -1230 669
rect -1331 634 -1298 668
rect -1264 634 -1230 668
rect -1974 566 -1940 600
rect -1906 566 -1873 600
rect -1974 532 -1873 566
rect -1974 498 -1940 532
rect -1906 498 -1873 532
rect -1974 298 -1873 498
rect -1974 264 -1940 298
rect -1906 264 -1873 298
rect -1974 230 -1873 264
rect -1974 196 -1940 230
rect -1906 196 -1873 230
rect -1974 162 -1873 196
rect -1811 583 -1393 607
rect -1811 549 -1787 583
rect -1753 549 -1719 583
rect -1685 549 -1519 583
rect -1485 549 -1451 583
rect -1417 549 -1393 583
rect -1811 535 -1393 549
rect -1811 515 -1739 535
rect -1811 481 -1787 515
rect -1753 481 -1739 515
rect -1811 315 -1739 481
rect -1465 515 -1393 535
rect -1465 481 -1451 515
rect -1417 481 -1393 515
rect -1681 463 -1523 477
rect -1681 429 -1667 463
rect -1633 449 -1571 463
rect -1537 429 -1523 463
rect -1681 367 -1653 429
rect -1551 367 -1523 429
rect -1681 333 -1667 367
rect -1633 333 -1571 347
rect -1537 333 -1523 367
rect -1681 319 -1523 333
rect -1811 281 -1787 315
rect -1753 281 -1739 315
rect -1811 261 -1739 281
rect -1465 315 -1393 481
rect -1465 281 -1451 315
rect -1417 281 -1393 315
rect -1465 261 -1393 281
rect -1811 247 -1393 261
rect -1811 213 -1787 247
rect -1753 213 -1719 247
rect -1685 213 -1519 247
rect -1485 213 -1451 247
rect -1417 213 -1393 247
rect -1811 189 -1393 213
rect -1331 600 -1230 634
rect -1331 566 -1298 600
rect -1264 566 -1230 600
rect -1331 532 -1230 566
rect -1331 498 -1298 532
rect -1264 498 -1230 532
rect -1331 298 -1230 498
rect -1331 264 -1298 298
rect -1264 264 -1230 298
rect -1331 230 -1230 264
rect -1331 196 -1298 230
rect -1264 196 -1230 230
rect -1974 128 -1940 162
rect -1906 128 -1873 162
rect -1974 127 -1873 128
rect -1331 162 -1230 196
rect -1331 128 -1298 162
rect -1264 128 -1230 162
rect -1331 127 -1230 128
rect -1974 94 -1230 127
rect -1974 60 -1940 94
rect -1906 60 -1872 94
rect -1838 60 -1804 94
rect -1770 60 -1736 94
rect -1702 60 -1502 94
rect -1468 60 -1434 94
rect -1400 60 -1366 94
rect -1332 60 -1298 94
rect -1264 60 -1230 94
rect -1974 26 -1230 60
rect -974 736 -230 770
rect -974 702 -940 736
rect -906 702 -872 736
rect -838 702 -804 736
rect -770 702 -736 736
rect -702 702 -502 736
rect -468 702 -434 736
rect -400 702 -366 736
rect -332 702 -298 736
rect -264 702 -230 736
rect -974 669 -230 702
rect -974 668 -873 669
rect -974 634 -940 668
rect -906 634 -873 668
rect -974 600 -873 634
rect -331 668 -230 669
rect -331 634 -298 668
rect -264 634 -230 668
rect -974 566 -940 600
rect -906 566 -873 600
rect -974 532 -873 566
rect -974 498 -940 532
rect -906 498 -873 532
rect -974 298 -873 498
rect -974 264 -940 298
rect -906 264 -873 298
rect -974 230 -873 264
rect -974 196 -940 230
rect -906 196 -873 230
rect -974 162 -873 196
rect -811 583 -393 607
rect -811 549 -787 583
rect -753 549 -719 583
rect -685 549 -519 583
rect -485 549 -451 583
rect -417 549 -393 583
rect -811 535 -393 549
rect -811 515 -739 535
rect -811 481 -787 515
rect -753 481 -739 515
rect -811 315 -739 481
rect -465 515 -393 535
rect -465 481 -451 515
rect -417 481 -393 515
rect -681 463 -523 477
rect -681 429 -667 463
rect -633 449 -571 463
rect -537 429 -523 463
rect -681 367 -653 429
rect -551 367 -523 429
rect -681 333 -667 367
rect -633 333 -571 347
rect -537 333 -523 367
rect -681 319 -523 333
rect -811 281 -787 315
rect -753 281 -739 315
rect -811 261 -739 281
rect -465 315 -393 481
rect -465 281 -451 315
rect -417 281 -393 315
rect -465 261 -393 281
rect -811 247 -393 261
rect -811 213 -787 247
rect -753 213 -719 247
rect -685 213 -519 247
rect -485 213 -451 247
rect -417 213 -393 247
rect -811 189 -393 213
rect -331 600 -230 634
rect -331 566 -298 600
rect -264 566 -230 600
rect -331 532 -230 566
rect -331 498 -298 532
rect -264 498 -230 532
rect -331 298 -230 498
rect -331 264 -298 298
rect -264 264 -230 298
rect -331 230 -230 264
rect -331 196 -298 230
rect -264 196 -230 230
rect -974 128 -940 162
rect -906 128 -873 162
rect -974 127 -873 128
rect -331 162 -230 196
rect -331 128 -298 162
rect -264 128 -230 162
rect -331 127 -230 128
rect -974 94 -230 127
rect -974 60 -940 94
rect -906 60 -872 94
rect -838 60 -804 94
rect -770 60 -736 94
rect -702 60 -502 94
rect -468 60 -434 94
rect -400 60 -366 94
rect -332 60 -298 94
rect -264 60 -230 94
rect -974 26 -230 60
rect 1026 736 1770 770
rect 1026 702 1060 736
rect 1094 702 1128 736
rect 1162 702 1196 736
rect 1230 702 1264 736
rect 1298 702 1498 736
rect 1532 702 1566 736
rect 1600 702 1634 736
rect 1668 702 1702 736
rect 1736 702 1770 736
rect 1026 669 1770 702
rect 1026 668 1127 669
rect 1026 634 1060 668
rect 1094 634 1127 668
rect 1026 600 1127 634
rect 1669 668 1770 669
rect 1669 634 1702 668
rect 1736 634 1770 668
rect 1026 566 1060 600
rect 1094 566 1127 600
rect 1026 532 1127 566
rect 1026 498 1060 532
rect 1094 498 1127 532
rect 1026 298 1127 498
rect 1026 264 1060 298
rect 1094 264 1127 298
rect 1026 230 1127 264
rect 1026 196 1060 230
rect 1094 196 1127 230
rect 1026 162 1127 196
rect 1189 583 1607 607
rect 1189 549 1213 583
rect 1247 549 1281 583
rect 1315 549 1481 583
rect 1515 549 1549 583
rect 1583 549 1607 583
rect 1189 535 1607 549
rect 1189 515 1261 535
rect 1189 481 1213 515
rect 1247 481 1261 515
rect 1189 315 1261 481
rect 1535 515 1607 535
rect 1535 481 1549 515
rect 1583 481 1607 515
rect 1319 463 1477 477
rect 1319 429 1333 463
rect 1367 449 1429 463
rect 1463 429 1477 463
rect 1319 367 1347 429
rect 1449 367 1477 429
rect 1319 333 1333 367
rect 1367 333 1429 347
rect 1463 333 1477 367
rect 1319 319 1477 333
rect 1189 281 1213 315
rect 1247 281 1261 315
rect 1189 261 1261 281
rect 1535 315 1607 481
rect 1535 281 1549 315
rect 1583 281 1607 315
rect 1535 261 1607 281
rect 1189 247 1607 261
rect 1189 213 1213 247
rect 1247 213 1281 247
rect 1315 213 1481 247
rect 1515 213 1549 247
rect 1583 213 1607 247
rect 1189 189 1607 213
rect 1669 600 1770 634
rect 1669 566 1702 600
rect 1736 566 1770 600
rect 1669 532 1770 566
rect 1669 498 1702 532
rect 1736 498 1770 532
rect 1669 298 1770 498
rect 1669 264 1702 298
rect 1736 264 1770 298
rect 1669 230 1770 264
rect 1669 196 1702 230
rect 1736 196 1770 230
rect 1026 128 1060 162
rect 1094 128 1127 162
rect 1026 127 1127 128
rect 1669 162 1770 196
rect 1669 128 1702 162
rect 1736 128 1770 162
rect 1669 127 1770 128
rect 1026 94 1770 127
rect 1026 60 1060 94
rect 1094 60 1128 94
rect 1162 60 1196 94
rect 1230 60 1264 94
rect 1298 60 1498 94
rect 1532 60 1566 94
rect 1600 60 1634 94
rect 1668 60 1702 94
rect 1736 60 1770 94
rect 1026 26 1770 60
rect 2026 736 2770 770
rect 2026 702 2060 736
rect 2094 702 2128 736
rect 2162 702 2196 736
rect 2230 702 2264 736
rect 2298 702 2498 736
rect 2532 702 2566 736
rect 2600 702 2634 736
rect 2668 702 2702 736
rect 2736 702 2770 736
rect 2026 669 2770 702
rect 2026 668 2127 669
rect 2026 634 2060 668
rect 2094 634 2127 668
rect 2026 600 2127 634
rect 2669 668 2770 669
rect 2669 634 2702 668
rect 2736 634 2770 668
rect 2026 566 2060 600
rect 2094 566 2127 600
rect 2026 532 2127 566
rect 2026 498 2060 532
rect 2094 498 2127 532
rect 2026 298 2127 498
rect 2026 264 2060 298
rect 2094 264 2127 298
rect 2026 230 2127 264
rect 2026 196 2060 230
rect 2094 196 2127 230
rect 2026 162 2127 196
rect 2189 583 2607 607
rect 2189 549 2213 583
rect 2247 549 2281 583
rect 2315 549 2481 583
rect 2515 549 2549 583
rect 2583 549 2607 583
rect 2189 535 2607 549
rect 2189 515 2261 535
rect 2189 481 2213 515
rect 2247 481 2261 515
rect 2189 315 2261 481
rect 2535 515 2607 535
rect 2535 481 2549 515
rect 2583 481 2607 515
rect 2319 463 2477 477
rect 2319 429 2333 463
rect 2367 449 2429 463
rect 2463 429 2477 463
rect 2319 367 2347 429
rect 2449 367 2477 429
rect 2319 333 2333 367
rect 2367 333 2429 347
rect 2463 333 2477 367
rect 2319 319 2477 333
rect 2189 281 2213 315
rect 2247 281 2261 315
rect 2189 261 2261 281
rect 2535 315 2607 481
rect 2535 281 2549 315
rect 2583 281 2607 315
rect 2535 261 2607 281
rect 2189 247 2607 261
rect 2189 213 2213 247
rect 2247 213 2281 247
rect 2315 213 2481 247
rect 2515 213 2549 247
rect 2583 213 2607 247
rect 2189 189 2607 213
rect 2669 600 2770 634
rect 2669 566 2702 600
rect 2736 566 2770 600
rect 2669 532 2770 566
rect 2669 498 2702 532
rect 2736 498 2770 532
rect 2669 298 2770 498
rect 2669 264 2702 298
rect 2736 264 2770 298
rect 2669 230 2770 264
rect 2669 196 2702 230
rect 2736 196 2770 230
rect 2026 128 2060 162
rect 2094 128 2127 162
rect 2026 127 2127 128
rect 2669 162 2770 196
rect 2669 128 2702 162
rect 2736 128 2770 162
rect 2669 127 2770 128
rect 2026 94 2770 127
rect 2026 60 2060 94
rect 2094 60 2128 94
rect 2162 60 2196 94
rect 2230 60 2264 94
rect 2298 60 2498 94
rect 2532 60 2566 94
rect 2600 60 2634 94
rect 2668 60 2702 94
rect 2736 60 2770 94
rect 2026 26 2770 60
rect 3026 736 3770 770
rect 3026 702 3060 736
rect 3094 702 3128 736
rect 3162 702 3196 736
rect 3230 702 3264 736
rect 3298 702 3498 736
rect 3532 702 3566 736
rect 3600 702 3634 736
rect 3668 702 3702 736
rect 3736 702 3770 736
rect 3026 669 3770 702
rect 3026 668 3127 669
rect 3026 634 3060 668
rect 3094 634 3127 668
rect 3026 600 3127 634
rect 3669 668 3770 669
rect 3669 634 3702 668
rect 3736 634 3770 668
rect 3026 566 3060 600
rect 3094 566 3127 600
rect 3026 532 3127 566
rect 3026 498 3060 532
rect 3094 498 3127 532
rect 3026 298 3127 498
rect 3026 264 3060 298
rect 3094 264 3127 298
rect 3026 230 3127 264
rect 3026 196 3060 230
rect 3094 196 3127 230
rect 3026 162 3127 196
rect 3189 583 3607 607
rect 3189 549 3213 583
rect 3247 549 3281 583
rect 3315 549 3481 583
rect 3515 549 3549 583
rect 3583 549 3607 583
rect 3189 535 3607 549
rect 3189 515 3261 535
rect 3189 481 3213 515
rect 3247 481 3261 515
rect 3189 315 3261 481
rect 3535 515 3607 535
rect 3535 481 3549 515
rect 3583 481 3607 515
rect 3319 463 3477 477
rect 3319 429 3333 463
rect 3367 449 3429 463
rect 3463 429 3477 463
rect 3319 367 3347 429
rect 3449 367 3477 429
rect 3319 333 3333 367
rect 3367 333 3429 347
rect 3463 333 3477 367
rect 3319 319 3477 333
rect 3189 281 3213 315
rect 3247 281 3261 315
rect 3189 261 3261 281
rect 3535 315 3607 481
rect 3535 281 3549 315
rect 3583 281 3607 315
rect 3535 261 3607 281
rect 3189 247 3607 261
rect 3189 213 3213 247
rect 3247 213 3281 247
rect 3315 213 3481 247
rect 3515 213 3549 247
rect 3583 213 3607 247
rect 3189 189 3607 213
rect 3669 600 3770 634
rect 3669 566 3702 600
rect 3736 566 3770 600
rect 3669 532 3770 566
rect 3669 498 3702 532
rect 3736 498 3770 532
rect 3669 298 3770 498
rect 3669 264 3702 298
rect 3736 264 3770 298
rect 3669 230 3770 264
rect 3669 196 3702 230
rect 3736 196 3770 230
rect 3026 128 3060 162
rect 3094 128 3127 162
rect 3026 127 3127 128
rect 3669 162 3770 196
rect 3669 128 3702 162
rect 3736 128 3770 162
rect 3669 127 3770 128
rect 3026 94 3770 127
rect 3026 60 3060 94
rect 3094 60 3128 94
rect 3162 60 3196 94
rect 3230 60 3264 94
rect 3298 60 3498 94
rect 3532 60 3566 94
rect 3600 60 3634 94
rect 3668 60 3702 94
rect 3736 60 3770 94
rect 3026 26 3770 60
rect -3974 -264 -3230 -230
rect -3974 -298 -3940 -264
rect -3906 -298 -3872 -264
rect -3838 -298 -3804 -264
rect -3770 -298 -3736 -264
rect -3702 -298 -3502 -264
rect -3468 -298 -3434 -264
rect -3400 -298 -3366 -264
rect -3332 -298 -3298 -264
rect -3264 -298 -3230 -264
rect -3974 -331 -3230 -298
rect -3974 -332 -3873 -331
rect -3974 -366 -3940 -332
rect -3906 -366 -3873 -332
rect -3974 -400 -3873 -366
rect -3331 -332 -3230 -331
rect -3331 -366 -3298 -332
rect -3264 -366 -3230 -332
rect -3974 -434 -3940 -400
rect -3906 -434 -3873 -400
rect -3974 -468 -3873 -434
rect -3974 -502 -3940 -468
rect -3906 -502 -3873 -468
rect -3974 -702 -3873 -502
rect -3974 -736 -3940 -702
rect -3906 -736 -3873 -702
rect -3974 -770 -3873 -736
rect -3974 -804 -3940 -770
rect -3906 -804 -3873 -770
rect -3974 -838 -3873 -804
rect -3811 -417 -3393 -393
rect -3811 -451 -3787 -417
rect -3753 -451 -3719 -417
rect -3685 -451 -3519 -417
rect -3485 -451 -3451 -417
rect -3417 -451 -3393 -417
rect -3811 -465 -3393 -451
rect -3811 -485 -3739 -465
rect -3811 -519 -3787 -485
rect -3753 -519 -3739 -485
rect -3811 -685 -3739 -519
rect -3465 -485 -3393 -465
rect -3465 -519 -3451 -485
rect -3417 -519 -3393 -485
rect -3681 -537 -3523 -523
rect -3681 -571 -3667 -537
rect -3633 -551 -3571 -537
rect -3537 -571 -3523 -537
rect -3681 -633 -3653 -571
rect -3551 -633 -3523 -571
rect -3681 -667 -3667 -633
rect -3633 -667 -3571 -653
rect -3537 -667 -3523 -633
rect -3681 -681 -3523 -667
rect -3811 -719 -3787 -685
rect -3753 -719 -3739 -685
rect -3811 -739 -3739 -719
rect -3465 -685 -3393 -519
rect -3465 -719 -3451 -685
rect -3417 -719 -3393 -685
rect -3465 -739 -3393 -719
rect -3811 -753 -3393 -739
rect -3811 -787 -3787 -753
rect -3753 -787 -3719 -753
rect -3685 -787 -3519 -753
rect -3485 -787 -3451 -753
rect -3417 -787 -3393 -753
rect -3811 -811 -3393 -787
rect -3331 -400 -3230 -366
rect -3331 -434 -3298 -400
rect -3264 -434 -3230 -400
rect -3331 -468 -3230 -434
rect -3331 -502 -3298 -468
rect -3264 -502 -3230 -468
rect -3331 -702 -3230 -502
rect -3331 -736 -3298 -702
rect -3264 -736 -3230 -702
rect -3331 -770 -3230 -736
rect -3331 -804 -3298 -770
rect -3264 -804 -3230 -770
rect -3974 -872 -3940 -838
rect -3906 -872 -3873 -838
rect -3974 -873 -3873 -872
rect -3331 -838 -3230 -804
rect -3331 -872 -3298 -838
rect -3264 -872 -3230 -838
rect -3331 -873 -3230 -872
rect -3974 -906 -3230 -873
rect -3974 -940 -3940 -906
rect -3906 -940 -3872 -906
rect -3838 -940 -3804 -906
rect -3770 -940 -3736 -906
rect -3702 -940 -3502 -906
rect -3468 -940 -3434 -906
rect -3400 -940 -3366 -906
rect -3332 -940 -3298 -906
rect -3264 -940 -3230 -906
rect -3974 -974 -3230 -940
rect -2974 -264 -2230 -230
rect -2974 -298 -2940 -264
rect -2906 -298 -2872 -264
rect -2838 -298 -2804 -264
rect -2770 -298 -2736 -264
rect -2702 -298 -2502 -264
rect -2468 -298 -2434 -264
rect -2400 -298 -2366 -264
rect -2332 -298 -2298 -264
rect -2264 -298 -2230 -264
rect -2974 -331 -2230 -298
rect -2974 -332 -2873 -331
rect -2974 -366 -2940 -332
rect -2906 -366 -2873 -332
rect -2974 -400 -2873 -366
rect -2331 -332 -2230 -331
rect -2331 -366 -2298 -332
rect -2264 -366 -2230 -332
rect -2974 -434 -2940 -400
rect -2906 -434 -2873 -400
rect -2974 -468 -2873 -434
rect -2974 -502 -2940 -468
rect -2906 -502 -2873 -468
rect -2974 -702 -2873 -502
rect -2974 -736 -2940 -702
rect -2906 -736 -2873 -702
rect -2974 -770 -2873 -736
rect -2974 -804 -2940 -770
rect -2906 -804 -2873 -770
rect -2974 -838 -2873 -804
rect -2811 -417 -2393 -393
rect -2811 -451 -2787 -417
rect -2753 -451 -2719 -417
rect -2685 -451 -2519 -417
rect -2485 -451 -2451 -417
rect -2417 -451 -2393 -417
rect -2811 -465 -2393 -451
rect -2811 -485 -2739 -465
rect -2811 -519 -2787 -485
rect -2753 -519 -2739 -485
rect -2811 -685 -2739 -519
rect -2465 -485 -2393 -465
rect -2465 -519 -2451 -485
rect -2417 -519 -2393 -485
rect -2681 -537 -2523 -523
rect -2681 -571 -2667 -537
rect -2633 -551 -2571 -537
rect -2537 -571 -2523 -537
rect -2681 -633 -2653 -571
rect -2551 -633 -2523 -571
rect -2681 -667 -2667 -633
rect -2633 -667 -2571 -653
rect -2537 -667 -2523 -633
rect -2681 -681 -2523 -667
rect -2811 -719 -2787 -685
rect -2753 -719 -2739 -685
rect -2811 -739 -2739 -719
rect -2465 -685 -2393 -519
rect -2465 -719 -2451 -685
rect -2417 -719 -2393 -685
rect -2465 -739 -2393 -719
rect -2811 -753 -2393 -739
rect -2811 -787 -2787 -753
rect -2753 -787 -2719 -753
rect -2685 -787 -2519 -753
rect -2485 -787 -2451 -753
rect -2417 -787 -2393 -753
rect -2811 -811 -2393 -787
rect -2331 -400 -2230 -366
rect -2331 -434 -2298 -400
rect -2264 -434 -2230 -400
rect -2331 -468 -2230 -434
rect -2331 -502 -2298 -468
rect -2264 -502 -2230 -468
rect -2331 -702 -2230 -502
rect -2331 -736 -2298 -702
rect -2264 -736 -2230 -702
rect -2331 -770 -2230 -736
rect -2331 -804 -2298 -770
rect -2264 -804 -2230 -770
rect -2974 -872 -2940 -838
rect -2906 -872 -2873 -838
rect -2974 -873 -2873 -872
rect -2331 -838 -2230 -804
rect -2331 -872 -2298 -838
rect -2264 -872 -2230 -838
rect -2331 -873 -2230 -872
rect -2974 -906 -2230 -873
rect -2974 -940 -2940 -906
rect -2906 -940 -2872 -906
rect -2838 -940 -2804 -906
rect -2770 -940 -2736 -906
rect -2702 -940 -2502 -906
rect -2468 -940 -2434 -906
rect -2400 -940 -2366 -906
rect -2332 -940 -2298 -906
rect -2264 -940 -2230 -906
rect -2974 -974 -2230 -940
rect -1974 -264 -1230 -230
rect -1974 -298 -1940 -264
rect -1906 -298 -1872 -264
rect -1838 -298 -1804 -264
rect -1770 -298 -1736 -264
rect -1702 -298 -1502 -264
rect -1468 -298 -1434 -264
rect -1400 -298 -1366 -264
rect -1332 -298 -1298 -264
rect -1264 -298 -1230 -264
rect -1974 -331 -1230 -298
rect -1974 -332 -1873 -331
rect -1974 -366 -1940 -332
rect -1906 -366 -1873 -332
rect -1974 -400 -1873 -366
rect -1331 -332 -1230 -331
rect -1331 -366 -1298 -332
rect -1264 -366 -1230 -332
rect -1974 -434 -1940 -400
rect -1906 -434 -1873 -400
rect -1974 -468 -1873 -434
rect -1974 -502 -1940 -468
rect -1906 -502 -1873 -468
rect -1974 -702 -1873 -502
rect -1974 -736 -1940 -702
rect -1906 -736 -1873 -702
rect -1974 -770 -1873 -736
rect -1974 -804 -1940 -770
rect -1906 -804 -1873 -770
rect -1974 -838 -1873 -804
rect -1811 -417 -1393 -393
rect -1811 -451 -1787 -417
rect -1753 -451 -1719 -417
rect -1685 -451 -1519 -417
rect -1485 -451 -1451 -417
rect -1417 -451 -1393 -417
rect -1811 -465 -1393 -451
rect -1811 -485 -1739 -465
rect -1811 -519 -1787 -485
rect -1753 -519 -1739 -485
rect -1811 -685 -1739 -519
rect -1465 -485 -1393 -465
rect -1465 -519 -1451 -485
rect -1417 -519 -1393 -485
rect -1681 -537 -1523 -523
rect -1681 -571 -1667 -537
rect -1633 -551 -1571 -537
rect -1537 -571 -1523 -537
rect -1681 -633 -1653 -571
rect -1551 -633 -1523 -571
rect -1681 -667 -1667 -633
rect -1633 -667 -1571 -653
rect -1537 -667 -1523 -633
rect -1681 -681 -1523 -667
rect -1811 -719 -1787 -685
rect -1753 -719 -1739 -685
rect -1811 -739 -1739 -719
rect -1465 -685 -1393 -519
rect -1465 -719 -1451 -685
rect -1417 -719 -1393 -685
rect -1465 -739 -1393 -719
rect -1811 -753 -1393 -739
rect -1811 -787 -1787 -753
rect -1753 -787 -1719 -753
rect -1685 -787 -1519 -753
rect -1485 -787 -1451 -753
rect -1417 -787 -1393 -753
rect -1811 -811 -1393 -787
rect -1331 -400 -1230 -366
rect -1331 -434 -1298 -400
rect -1264 -434 -1230 -400
rect -1331 -468 -1230 -434
rect -1331 -502 -1298 -468
rect -1264 -502 -1230 -468
rect -1331 -702 -1230 -502
rect -1331 -736 -1298 -702
rect -1264 -736 -1230 -702
rect -1331 -770 -1230 -736
rect -1331 -804 -1298 -770
rect -1264 -804 -1230 -770
rect -1974 -872 -1940 -838
rect -1906 -872 -1873 -838
rect -1974 -873 -1873 -872
rect -1331 -838 -1230 -804
rect -1331 -872 -1298 -838
rect -1264 -872 -1230 -838
rect -1331 -873 -1230 -872
rect -1974 -906 -1230 -873
rect -1974 -940 -1940 -906
rect -1906 -940 -1872 -906
rect -1838 -940 -1804 -906
rect -1770 -940 -1736 -906
rect -1702 -940 -1502 -906
rect -1468 -940 -1434 -906
rect -1400 -940 -1366 -906
rect -1332 -940 -1298 -906
rect -1264 -940 -1230 -906
rect -1974 -974 -1230 -940
rect -974 -264 -230 -230
rect -974 -298 -940 -264
rect -906 -298 -872 -264
rect -838 -298 -804 -264
rect -770 -298 -736 -264
rect -702 -298 -502 -264
rect -468 -298 -434 -264
rect -400 -298 -366 -264
rect -332 -298 -298 -264
rect -264 -298 -230 -264
rect -974 -331 -230 -298
rect -974 -332 -873 -331
rect -974 -366 -940 -332
rect -906 -366 -873 -332
rect -974 -400 -873 -366
rect -331 -332 -230 -331
rect -331 -366 -298 -332
rect -264 -366 -230 -332
rect -974 -434 -940 -400
rect -906 -434 -873 -400
rect -974 -468 -873 -434
rect -974 -502 -940 -468
rect -906 -502 -873 -468
rect -974 -702 -873 -502
rect -974 -736 -940 -702
rect -906 -736 -873 -702
rect -974 -770 -873 -736
rect -974 -804 -940 -770
rect -906 -804 -873 -770
rect -974 -838 -873 -804
rect -811 -417 -393 -393
rect -811 -451 -787 -417
rect -753 -451 -719 -417
rect -685 -451 -519 -417
rect -485 -451 -451 -417
rect -417 -451 -393 -417
rect -811 -465 -393 -451
rect -811 -485 -739 -465
rect -811 -519 -787 -485
rect -753 -519 -739 -485
rect -811 -685 -739 -519
rect -465 -485 -393 -465
rect -465 -519 -451 -485
rect -417 -519 -393 -485
rect -681 -537 -523 -523
rect -681 -571 -667 -537
rect -633 -551 -571 -537
rect -537 -571 -523 -537
rect -681 -633 -653 -571
rect -551 -633 -523 -571
rect -681 -667 -667 -633
rect -633 -667 -571 -653
rect -537 -667 -523 -633
rect -681 -681 -523 -667
rect -811 -719 -787 -685
rect -753 -719 -739 -685
rect -811 -739 -739 -719
rect -465 -685 -393 -519
rect -465 -719 -451 -685
rect -417 -719 -393 -685
rect -465 -739 -393 -719
rect -811 -753 -393 -739
rect -811 -787 -787 -753
rect -753 -787 -719 -753
rect -685 -787 -519 -753
rect -485 -787 -451 -753
rect -417 -787 -393 -753
rect -811 -811 -393 -787
rect -331 -400 -230 -366
rect -331 -434 -298 -400
rect -264 -434 -230 -400
rect -331 -468 -230 -434
rect -331 -502 -298 -468
rect -264 -502 -230 -468
rect -331 -702 -230 -502
rect -331 -736 -298 -702
rect -264 -736 -230 -702
rect -331 -770 -230 -736
rect -331 -804 -298 -770
rect -264 -804 -230 -770
rect -974 -872 -940 -838
rect -906 -872 -873 -838
rect -974 -873 -873 -872
rect -331 -838 -230 -804
rect -331 -872 -298 -838
rect -264 -872 -230 -838
rect -331 -873 -230 -872
rect -974 -906 -230 -873
rect -974 -940 -940 -906
rect -906 -940 -872 -906
rect -838 -940 -804 -906
rect -770 -940 -736 -906
rect -702 -940 -502 -906
rect -468 -940 -434 -906
rect -400 -940 -366 -906
rect -332 -940 -298 -906
rect -264 -940 -230 -906
rect -974 -974 -230 -940
rect 26 -264 770 -230
rect 26 -298 60 -264
rect 94 -298 128 -264
rect 162 -298 196 -264
rect 230 -298 264 -264
rect 298 -298 498 -264
rect 532 -298 566 -264
rect 600 -298 634 -264
rect 668 -298 702 -264
rect 736 -298 770 -264
rect 26 -331 770 -298
rect 26 -332 127 -331
rect 26 -366 60 -332
rect 94 -366 127 -332
rect 26 -400 127 -366
rect 669 -332 770 -331
rect 669 -366 702 -332
rect 736 -366 770 -332
rect 26 -434 60 -400
rect 94 -434 127 -400
rect 26 -468 127 -434
rect 26 -502 60 -468
rect 94 -502 127 -468
rect 26 -702 127 -502
rect 26 -736 60 -702
rect 94 -736 127 -702
rect 26 -770 127 -736
rect 26 -804 60 -770
rect 94 -804 127 -770
rect 26 -838 127 -804
rect 189 -417 607 -393
rect 189 -451 213 -417
rect 247 -451 281 -417
rect 315 -451 481 -417
rect 515 -451 549 -417
rect 583 -451 607 -417
rect 189 -465 607 -451
rect 189 -485 261 -465
rect 189 -519 213 -485
rect 247 -519 261 -485
rect 189 -685 261 -519
rect 535 -485 607 -465
rect 535 -519 549 -485
rect 583 -519 607 -485
rect 319 -537 477 -523
rect 319 -571 333 -537
rect 367 -551 429 -537
rect 463 -571 477 -537
rect 319 -633 347 -571
rect 449 -633 477 -571
rect 319 -667 333 -633
rect 367 -667 429 -653
rect 463 -667 477 -633
rect 319 -681 477 -667
rect 189 -719 213 -685
rect 247 -719 261 -685
rect 189 -739 261 -719
rect 535 -685 607 -519
rect 535 -719 549 -685
rect 583 -719 607 -685
rect 535 -739 607 -719
rect 189 -753 607 -739
rect 189 -787 213 -753
rect 247 -787 281 -753
rect 315 -787 481 -753
rect 515 -787 549 -753
rect 583 -787 607 -753
rect 189 -811 607 -787
rect 669 -400 770 -366
rect 669 -434 702 -400
rect 736 -434 770 -400
rect 669 -468 770 -434
rect 669 -502 702 -468
rect 736 -502 770 -468
rect 669 -702 770 -502
rect 669 -736 702 -702
rect 736 -736 770 -702
rect 669 -770 770 -736
rect 669 -804 702 -770
rect 736 -804 770 -770
rect 26 -872 60 -838
rect 94 -872 127 -838
rect 26 -873 127 -872
rect 669 -838 770 -804
rect 669 -872 702 -838
rect 736 -872 770 -838
rect 669 -873 770 -872
rect 26 -906 770 -873
rect 26 -940 60 -906
rect 94 -940 128 -906
rect 162 -940 196 -906
rect 230 -940 264 -906
rect 298 -940 498 -906
rect 532 -940 566 -906
rect 600 -940 634 -906
rect 668 -940 702 -906
rect 736 -940 770 -906
rect 26 -974 770 -940
rect 1026 -264 1770 -230
rect 1026 -298 1060 -264
rect 1094 -298 1128 -264
rect 1162 -298 1196 -264
rect 1230 -298 1264 -264
rect 1298 -298 1498 -264
rect 1532 -298 1566 -264
rect 1600 -298 1634 -264
rect 1668 -298 1702 -264
rect 1736 -298 1770 -264
rect 1026 -331 1770 -298
rect 1026 -332 1127 -331
rect 1026 -366 1060 -332
rect 1094 -366 1127 -332
rect 1026 -400 1127 -366
rect 1669 -332 1770 -331
rect 1669 -366 1702 -332
rect 1736 -366 1770 -332
rect 1026 -434 1060 -400
rect 1094 -434 1127 -400
rect 1026 -468 1127 -434
rect 1026 -502 1060 -468
rect 1094 -502 1127 -468
rect 1026 -702 1127 -502
rect 1026 -736 1060 -702
rect 1094 -736 1127 -702
rect 1026 -770 1127 -736
rect 1026 -804 1060 -770
rect 1094 -804 1127 -770
rect 1026 -838 1127 -804
rect 1189 -417 1607 -393
rect 1189 -451 1213 -417
rect 1247 -451 1281 -417
rect 1315 -451 1481 -417
rect 1515 -451 1549 -417
rect 1583 -451 1607 -417
rect 1189 -465 1607 -451
rect 1189 -485 1261 -465
rect 1189 -519 1213 -485
rect 1247 -519 1261 -485
rect 1189 -685 1261 -519
rect 1535 -485 1607 -465
rect 1535 -519 1549 -485
rect 1583 -519 1607 -485
rect 1319 -537 1477 -523
rect 1319 -571 1333 -537
rect 1367 -551 1429 -537
rect 1463 -571 1477 -537
rect 1319 -633 1347 -571
rect 1449 -633 1477 -571
rect 1319 -667 1333 -633
rect 1367 -667 1429 -653
rect 1463 -667 1477 -633
rect 1319 -681 1477 -667
rect 1189 -719 1213 -685
rect 1247 -719 1261 -685
rect 1189 -739 1261 -719
rect 1535 -685 1607 -519
rect 1535 -719 1549 -685
rect 1583 -719 1607 -685
rect 1535 -739 1607 -719
rect 1189 -753 1607 -739
rect 1189 -787 1213 -753
rect 1247 -787 1281 -753
rect 1315 -787 1481 -753
rect 1515 -787 1549 -753
rect 1583 -787 1607 -753
rect 1189 -811 1607 -787
rect 1669 -400 1770 -366
rect 1669 -434 1702 -400
rect 1736 -434 1770 -400
rect 1669 -468 1770 -434
rect 1669 -502 1702 -468
rect 1736 -502 1770 -468
rect 1669 -702 1770 -502
rect 1669 -736 1702 -702
rect 1736 -736 1770 -702
rect 1669 -770 1770 -736
rect 1669 -804 1702 -770
rect 1736 -804 1770 -770
rect 1026 -872 1060 -838
rect 1094 -872 1127 -838
rect 1026 -873 1127 -872
rect 1669 -838 1770 -804
rect 1669 -872 1702 -838
rect 1736 -872 1770 -838
rect 1669 -873 1770 -872
rect 1026 -906 1770 -873
rect 1026 -940 1060 -906
rect 1094 -940 1128 -906
rect 1162 -940 1196 -906
rect 1230 -940 1264 -906
rect 1298 -940 1498 -906
rect 1532 -940 1566 -906
rect 1600 -940 1634 -906
rect 1668 -940 1702 -906
rect 1736 -940 1770 -906
rect 1026 -974 1770 -940
rect 2026 -264 2770 -230
rect 2026 -298 2060 -264
rect 2094 -298 2128 -264
rect 2162 -298 2196 -264
rect 2230 -298 2264 -264
rect 2298 -298 2498 -264
rect 2532 -298 2566 -264
rect 2600 -298 2634 -264
rect 2668 -298 2702 -264
rect 2736 -298 2770 -264
rect 2026 -331 2770 -298
rect 2026 -332 2127 -331
rect 2026 -366 2060 -332
rect 2094 -366 2127 -332
rect 2026 -400 2127 -366
rect 2669 -332 2770 -331
rect 2669 -366 2702 -332
rect 2736 -366 2770 -332
rect 2026 -434 2060 -400
rect 2094 -434 2127 -400
rect 2026 -468 2127 -434
rect 2026 -502 2060 -468
rect 2094 -502 2127 -468
rect 2026 -702 2127 -502
rect 2026 -736 2060 -702
rect 2094 -736 2127 -702
rect 2026 -770 2127 -736
rect 2026 -804 2060 -770
rect 2094 -804 2127 -770
rect 2026 -838 2127 -804
rect 2189 -417 2607 -393
rect 2189 -451 2213 -417
rect 2247 -451 2281 -417
rect 2315 -451 2481 -417
rect 2515 -451 2549 -417
rect 2583 -451 2607 -417
rect 2189 -465 2607 -451
rect 2189 -485 2261 -465
rect 2189 -519 2213 -485
rect 2247 -519 2261 -485
rect 2189 -685 2261 -519
rect 2535 -485 2607 -465
rect 2535 -519 2549 -485
rect 2583 -519 2607 -485
rect 2319 -537 2477 -523
rect 2319 -571 2333 -537
rect 2367 -551 2429 -537
rect 2463 -571 2477 -537
rect 2319 -633 2347 -571
rect 2449 -633 2477 -571
rect 2319 -667 2333 -633
rect 2367 -667 2429 -653
rect 2463 -667 2477 -633
rect 2319 -681 2477 -667
rect 2189 -719 2213 -685
rect 2247 -719 2261 -685
rect 2189 -739 2261 -719
rect 2535 -685 2607 -519
rect 2535 -719 2549 -685
rect 2583 -719 2607 -685
rect 2535 -739 2607 -719
rect 2189 -753 2607 -739
rect 2189 -787 2213 -753
rect 2247 -787 2281 -753
rect 2315 -787 2481 -753
rect 2515 -787 2549 -753
rect 2583 -787 2607 -753
rect 2189 -811 2607 -787
rect 2669 -400 2770 -366
rect 2669 -434 2702 -400
rect 2736 -434 2770 -400
rect 2669 -468 2770 -434
rect 2669 -502 2702 -468
rect 2736 -502 2770 -468
rect 2669 -702 2770 -502
rect 2669 -736 2702 -702
rect 2736 -736 2770 -702
rect 2669 -770 2770 -736
rect 2669 -804 2702 -770
rect 2736 -804 2770 -770
rect 2026 -872 2060 -838
rect 2094 -872 2127 -838
rect 2026 -873 2127 -872
rect 2669 -838 2770 -804
rect 2669 -872 2702 -838
rect 2736 -872 2770 -838
rect 2669 -873 2770 -872
rect 2026 -906 2770 -873
rect 2026 -940 2060 -906
rect 2094 -940 2128 -906
rect 2162 -940 2196 -906
rect 2230 -940 2264 -906
rect 2298 -940 2498 -906
rect 2532 -940 2566 -906
rect 2600 -940 2634 -906
rect 2668 -940 2702 -906
rect 2736 -940 2770 -906
rect 2026 -974 2770 -940
rect 3026 -264 3770 -230
rect 3026 -298 3060 -264
rect 3094 -298 3128 -264
rect 3162 -298 3196 -264
rect 3230 -298 3264 -264
rect 3298 -298 3498 -264
rect 3532 -298 3566 -264
rect 3600 -298 3634 -264
rect 3668 -298 3702 -264
rect 3736 -298 3770 -264
rect 3026 -331 3770 -298
rect 3026 -332 3127 -331
rect 3026 -366 3060 -332
rect 3094 -366 3127 -332
rect 3026 -400 3127 -366
rect 3669 -332 3770 -331
rect 3669 -366 3702 -332
rect 3736 -366 3770 -332
rect 3026 -434 3060 -400
rect 3094 -434 3127 -400
rect 3026 -468 3127 -434
rect 3026 -502 3060 -468
rect 3094 -502 3127 -468
rect 3026 -702 3127 -502
rect 3026 -736 3060 -702
rect 3094 -736 3127 -702
rect 3026 -770 3127 -736
rect 3026 -804 3060 -770
rect 3094 -804 3127 -770
rect 3026 -838 3127 -804
rect 3189 -417 3607 -393
rect 3189 -451 3213 -417
rect 3247 -451 3281 -417
rect 3315 -451 3481 -417
rect 3515 -451 3549 -417
rect 3583 -451 3607 -417
rect 3189 -465 3607 -451
rect 3189 -485 3261 -465
rect 3189 -519 3213 -485
rect 3247 -519 3261 -485
rect 3189 -685 3261 -519
rect 3535 -485 3607 -465
rect 3535 -519 3549 -485
rect 3583 -519 3607 -485
rect 3319 -537 3477 -523
rect 3319 -571 3333 -537
rect 3367 -551 3429 -537
rect 3463 -571 3477 -537
rect 3319 -633 3347 -571
rect 3449 -633 3477 -571
rect 3319 -667 3333 -633
rect 3367 -667 3429 -653
rect 3463 -667 3477 -633
rect 3319 -681 3477 -667
rect 3189 -719 3213 -685
rect 3247 -719 3261 -685
rect 3189 -739 3261 -719
rect 3535 -685 3607 -519
rect 3535 -719 3549 -685
rect 3583 -719 3607 -685
rect 3535 -739 3607 -719
rect 3189 -753 3607 -739
rect 3189 -787 3213 -753
rect 3247 -787 3281 -753
rect 3315 -787 3481 -753
rect 3515 -787 3549 -753
rect 3583 -787 3607 -753
rect 3189 -811 3607 -787
rect 3669 -400 3770 -366
rect 3669 -434 3702 -400
rect 3736 -434 3770 -400
rect 3669 -468 3770 -434
rect 3669 -502 3702 -468
rect 3736 -502 3770 -468
rect 3669 -702 3770 -502
rect 3669 -736 3702 -702
rect 3736 -736 3770 -702
rect 3669 -770 3770 -736
rect 3669 -804 3702 -770
rect 3736 -804 3770 -770
rect 3026 -872 3060 -838
rect 3094 -872 3127 -838
rect 3026 -873 3127 -872
rect 3669 -838 3770 -804
rect 3669 -872 3702 -838
rect 3736 -872 3770 -838
rect 3669 -873 3770 -872
rect 3026 -906 3770 -873
rect 3026 -940 3060 -906
rect 3094 -940 3128 -906
rect 3162 -940 3196 -906
rect 3230 -940 3264 -906
rect 3298 -940 3498 -906
rect 3532 -940 3566 -906
rect 3600 -940 3634 -906
rect 3668 -940 3702 -906
rect 3736 -940 3770 -906
rect 3026 -974 3770 -940
rect -974 -1264 -230 -1230
rect -974 -1298 -940 -1264
rect -906 -1298 -872 -1264
rect -838 -1298 -804 -1264
rect -770 -1298 -736 -1264
rect -702 -1298 -502 -1264
rect -468 -1298 -434 -1264
rect -400 -1298 -366 -1264
rect -332 -1298 -298 -1264
rect -264 -1298 -230 -1264
rect -974 -1331 -230 -1298
rect -974 -1332 -873 -1331
rect -974 -1366 -940 -1332
rect -906 -1366 -873 -1332
rect -974 -1400 -873 -1366
rect -331 -1332 -230 -1331
rect -331 -1366 -298 -1332
rect -264 -1366 -230 -1332
rect -974 -1434 -940 -1400
rect -906 -1434 -873 -1400
rect -974 -1468 -873 -1434
rect -974 -1502 -940 -1468
rect -906 -1502 -873 -1468
rect -974 -1702 -873 -1502
rect -974 -1736 -940 -1702
rect -906 -1736 -873 -1702
rect -974 -1770 -873 -1736
rect -974 -1804 -940 -1770
rect -906 -1804 -873 -1770
rect -974 -1838 -873 -1804
rect -811 -1417 -393 -1393
rect -811 -1451 -787 -1417
rect -753 -1451 -719 -1417
rect -685 -1451 -519 -1417
rect -485 -1451 -451 -1417
rect -417 -1451 -393 -1417
rect -811 -1465 -393 -1451
rect -811 -1485 -739 -1465
rect -811 -1519 -787 -1485
rect -753 -1519 -739 -1485
rect -811 -1685 -739 -1519
rect -465 -1485 -393 -1465
rect -465 -1519 -451 -1485
rect -417 -1519 -393 -1485
rect -681 -1537 -523 -1523
rect -681 -1571 -667 -1537
rect -633 -1551 -571 -1537
rect -537 -1571 -523 -1537
rect -681 -1633 -653 -1571
rect -551 -1633 -523 -1571
rect -681 -1667 -667 -1633
rect -633 -1667 -571 -1653
rect -537 -1667 -523 -1633
rect -681 -1681 -523 -1667
rect -811 -1719 -787 -1685
rect -753 -1719 -739 -1685
rect -811 -1739 -739 -1719
rect -465 -1685 -393 -1519
rect -465 -1719 -451 -1685
rect -417 -1719 -393 -1685
rect -465 -1739 -393 -1719
rect -811 -1753 -393 -1739
rect -811 -1787 -787 -1753
rect -753 -1787 -719 -1753
rect -685 -1787 -519 -1753
rect -485 -1787 -451 -1753
rect -417 -1787 -393 -1753
rect -811 -1811 -393 -1787
rect -331 -1400 -230 -1366
rect -331 -1434 -298 -1400
rect -264 -1434 -230 -1400
rect -331 -1468 -230 -1434
rect -331 -1502 -298 -1468
rect -264 -1502 -230 -1468
rect -331 -1702 -230 -1502
rect -331 -1736 -298 -1702
rect -264 -1736 -230 -1702
rect -331 -1770 -230 -1736
rect -331 -1804 -298 -1770
rect -264 -1804 -230 -1770
rect -974 -1872 -940 -1838
rect -906 -1872 -873 -1838
rect -974 -1873 -873 -1872
rect -331 -1838 -230 -1804
rect -331 -1872 -298 -1838
rect -264 -1872 -230 -1838
rect -331 -1873 -230 -1872
rect -974 -1906 -230 -1873
rect -974 -1940 -940 -1906
rect -906 -1940 -872 -1906
rect -838 -1940 -804 -1906
rect -770 -1940 -736 -1906
rect -702 -1940 -502 -1906
rect -468 -1940 -434 -1906
rect -400 -1940 -366 -1906
rect -332 -1940 -298 -1906
rect -264 -1940 -230 -1906
rect -974 -1974 -230 -1940
rect 26 -1264 770 -1230
rect 26 -1298 60 -1264
rect 94 -1298 128 -1264
rect 162 -1298 196 -1264
rect 230 -1298 264 -1264
rect 298 -1298 498 -1264
rect 532 -1298 566 -1264
rect 600 -1298 634 -1264
rect 668 -1298 702 -1264
rect 736 -1298 770 -1264
rect 26 -1331 770 -1298
rect 26 -1332 127 -1331
rect 26 -1366 60 -1332
rect 94 -1366 127 -1332
rect 26 -1400 127 -1366
rect 669 -1332 770 -1331
rect 669 -1366 702 -1332
rect 736 -1366 770 -1332
rect 26 -1434 60 -1400
rect 94 -1434 127 -1400
rect 26 -1468 127 -1434
rect 26 -1502 60 -1468
rect 94 -1502 127 -1468
rect 26 -1702 127 -1502
rect 26 -1736 60 -1702
rect 94 -1736 127 -1702
rect 26 -1770 127 -1736
rect 26 -1804 60 -1770
rect 94 -1804 127 -1770
rect 26 -1838 127 -1804
rect 189 -1417 607 -1393
rect 189 -1451 213 -1417
rect 247 -1451 281 -1417
rect 315 -1451 481 -1417
rect 515 -1451 549 -1417
rect 583 -1451 607 -1417
rect 189 -1465 607 -1451
rect 189 -1485 261 -1465
rect 189 -1519 213 -1485
rect 247 -1519 261 -1485
rect 189 -1685 261 -1519
rect 535 -1485 607 -1465
rect 535 -1519 549 -1485
rect 583 -1519 607 -1485
rect 319 -1537 477 -1523
rect 319 -1571 333 -1537
rect 367 -1551 429 -1537
rect 463 -1571 477 -1537
rect 319 -1633 347 -1571
rect 449 -1633 477 -1571
rect 319 -1667 333 -1633
rect 367 -1667 429 -1653
rect 463 -1667 477 -1633
rect 319 -1681 477 -1667
rect 189 -1719 213 -1685
rect 247 -1719 261 -1685
rect 189 -1739 261 -1719
rect 535 -1685 607 -1519
rect 535 -1719 549 -1685
rect 583 -1719 607 -1685
rect 535 -1739 607 -1719
rect 189 -1753 607 -1739
rect 189 -1787 213 -1753
rect 247 -1787 281 -1753
rect 315 -1787 481 -1753
rect 515 -1787 549 -1753
rect 583 -1787 607 -1753
rect 189 -1811 607 -1787
rect 669 -1400 770 -1366
rect 669 -1434 702 -1400
rect 736 -1434 770 -1400
rect 669 -1468 770 -1434
rect 669 -1502 702 -1468
rect 736 -1502 770 -1468
rect 669 -1702 770 -1502
rect 669 -1736 702 -1702
rect 736 -1736 770 -1702
rect 669 -1770 770 -1736
rect 669 -1804 702 -1770
rect 736 -1804 770 -1770
rect 26 -1872 60 -1838
rect 94 -1872 127 -1838
rect 26 -1873 127 -1872
rect 669 -1838 770 -1804
rect 669 -1872 702 -1838
rect 736 -1872 770 -1838
rect 669 -1873 770 -1872
rect 26 -1906 770 -1873
rect 26 -1940 60 -1906
rect 94 -1940 128 -1906
rect 162 -1940 196 -1906
rect 230 -1940 264 -1906
rect 298 -1940 498 -1906
rect 532 -1940 566 -1906
rect 600 -1940 634 -1906
rect 668 -1940 702 -1906
rect 736 -1940 770 -1906
rect 26 -1974 770 -1940
rect 1026 -1264 1770 -1230
rect 1026 -1298 1060 -1264
rect 1094 -1298 1128 -1264
rect 1162 -1298 1196 -1264
rect 1230 -1298 1264 -1264
rect 1298 -1298 1498 -1264
rect 1532 -1298 1566 -1264
rect 1600 -1298 1634 -1264
rect 1668 -1298 1702 -1264
rect 1736 -1298 1770 -1264
rect 1026 -1331 1770 -1298
rect 1026 -1332 1127 -1331
rect 1026 -1366 1060 -1332
rect 1094 -1366 1127 -1332
rect 1026 -1400 1127 -1366
rect 1669 -1332 1770 -1331
rect 1669 -1366 1702 -1332
rect 1736 -1366 1770 -1332
rect 1026 -1434 1060 -1400
rect 1094 -1434 1127 -1400
rect 1026 -1468 1127 -1434
rect 1026 -1502 1060 -1468
rect 1094 -1502 1127 -1468
rect 1026 -1702 1127 -1502
rect 1026 -1736 1060 -1702
rect 1094 -1736 1127 -1702
rect 1026 -1770 1127 -1736
rect 1026 -1804 1060 -1770
rect 1094 -1804 1127 -1770
rect 1026 -1838 1127 -1804
rect 1189 -1417 1607 -1393
rect 1189 -1451 1213 -1417
rect 1247 -1451 1281 -1417
rect 1315 -1451 1481 -1417
rect 1515 -1451 1549 -1417
rect 1583 -1451 1607 -1417
rect 1189 -1465 1607 -1451
rect 1189 -1485 1261 -1465
rect 1189 -1519 1213 -1485
rect 1247 -1519 1261 -1485
rect 1189 -1685 1261 -1519
rect 1535 -1485 1607 -1465
rect 1535 -1519 1549 -1485
rect 1583 -1519 1607 -1485
rect 1319 -1537 1477 -1523
rect 1319 -1571 1333 -1537
rect 1367 -1551 1429 -1537
rect 1463 -1571 1477 -1537
rect 1319 -1633 1347 -1571
rect 1449 -1633 1477 -1571
rect 1319 -1667 1333 -1633
rect 1367 -1667 1429 -1653
rect 1463 -1667 1477 -1633
rect 1319 -1681 1477 -1667
rect 1189 -1719 1213 -1685
rect 1247 -1719 1261 -1685
rect 1189 -1739 1261 -1719
rect 1535 -1685 1607 -1519
rect 1535 -1719 1549 -1685
rect 1583 -1719 1607 -1685
rect 1535 -1739 1607 -1719
rect 1189 -1753 1607 -1739
rect 1189 -1787 1213 -1753
rect 1247 -1787 1281 -1753
rect 1315 -1787 1481 -1753
rect 1515 -1787 1549 -1753
rect 1583 -1787 1607 -1753
rect 1189 -1811 1607 -1787
rect 1669 -1400 1770 -1366
rect 1669 -1434 1702 -1400
rect 1736 -1434 1770 -1400
rect 1669 -1468 1770 -1434
rect 1669 -1502 1702 -1468
rect 1736 -1502 1770 -1468
rect 1669 -1702 1770 -1502
rect 1669 -1736 1702 -1702
rect 1736 -1736 1770 -1702
rect 1669 -1770 1770 -1736
rect 1669 -1804 1702 -1770
rect 1736 -1804 1770 -1770
rect 1026 -1872 1060 -1838
rect 1094 -1872 1127 -1838
rect 1026 -1873 1127 -1872
rect 1669 -1838 1770 -1804
rect 1669 -1872 1702 -1838
rect 1736 -1872 1770 -1838
rect 1669 -1873 1770 -1872
rect 1026 -1906 1770 -1873
rect 1026 -1940 1060 -1906
rect 1094 -1940 1128 -1906
rect 1162 -1940 1196 -1906
rect 1230 -1940 1264 -1906
rect 1298 -1940 1498 -1906
rect 1532 -1940 1566 -1906
rect 1600 -1940 1634 -1906
rect 1668 -1940 1702 -1906
rect 1736 -1940 1770 -1906
rect 1026 -1974 1770 -1940
rect 2026 -1264 2770 -1230
rect 2026 -1298 2060 -1264
rect 2094 -1298 2128 -1264
rect 2162 -1298 2196 -1264
rect 2230 -1298 2264 -1264
rect 2298 -1298 2498 -1264
rect 2532 -1298 2566 -1264
rect 2600 -1298 2634 -1264
rect 2668 -1298 2702 -1264
rect 2736 -1298 2770 -1264
rect 2026 -1331 2770 -1298
rect 2026 -1332 2127 -1331
rect 2026 -1366 2060 -1332
rect 2094 -1366 2127 -1332
rect 2026 -1400 2127 -1366
rect 2669 -1332 2770 -1331
rect 2669 -1366 2702 -1332
rect 2736 -1366 2770 -1332
rect 2026 -1434 2060 -1400
rect 2094 -1434 2127 -1400
rect 2026 -1468 2127 -1434
rect 2026 -1502 2060 -1468
rect 2094 -1502 2127 -1468
rect 2026 -1702 2127 -1502
rect 2026 -1736 2060 -1702
rect 2094 -1736 2127 -1702
rect 2026 -1770 2127 -1736
rect 2026 -1804 2060 -1770
rect 2094 -1804 2127 -1770
rect 2026 -1838 2127 -1804
rect 2189 -1417 2607 -1393
rect 2189 -1451 2213 -1417
rect 2247 -1451 2281 -1417
rect 2315 -1451 2481 -1417
rect 2515 -1451 2549 -1417
rect 2583 -1451 2607 -1417
rect 2189 -1465 2607 -1451
rect 2189 -1485 2261 -1465
rect 2189 -1519 2213 -1485
rect 2247 -1519 2261 -1485
rect 2189 -1685 2261 -1519
rect 2535 -1485 2607 -1465
rect 2535 -1519 2549 -1485
rect 2583 -1519 2607 -1485
rect 2319 -1537 2477 -1523
rect 2319 -1571 2333 -1537
rect 2367 -1551 2429 -1537
rect 2463 -1571 2477 -1537
rect 2319 -1633 2347 -1571
rect 2449 -1633 2477 -1571
rect 2319 -1667 2333 -1633
rect 2367 -1667 2429 -1653
rect 2463 -1667 2477 -1633
rect 2319 -1681 2477 -1667
rect 2189 -1719 2213 -1685
rect 2247 -1719 2261 -1685
rect 2189 -1739 2261 -1719
rect 2535 -1685 2607 -1519
rect 2535 -1719 2549 -1685
rect 2583 -1719 2607 -1685
rect 2535 -1739 2607 -1719
rect 2189 -1753 2607 -1739
rect 2189 -1787 2213 -1753
rect 2247 -1787 2281 -1753
rect 2315 -1787 2481 -1753
rect 2515 -1787 2549 -1753
rect 2583 -1787 2607 -1753
rect 2189 -1811 2607 -1787
rect 2669 -1400 2770 -1366
rect 2669 -1434 2702 -1400
rect 2736 -1434 2770 -1400
rect 2669 -1468 2770 -1434
rect 2669 -1502 2702 -1468
rect 2736 -1502 2770 -1468
rect 2669 -1702 2770 -1502
rect 2669 -1736 2702 -1702
rect 2736 -1736 2770 -1702
rect 2669 -1770 2770 -1736
rect 2669 -1804 2702 -1770
rect 2736 -1804 2770 -1770
rect 2026 -1872 2060 -1838
rect 2094 -1872 2127 -1838
rect 2026 -1873 2127 -1872
rect 2669 -1838 2770 -1804
rect 2669 -1872 2702 -1838
rect 2736 -1872 2770 -1838
rect 2669 -1873 2770 -1872
rect 2026 -1906 2770 -1873
rect 2026 -1940 2060 -1906
rect 2094 -1940 2128 -1906
rect 2162 -1940 2196 -1906
rect 2230 -1940 2264 -1906
rect 2298 -1940 2498 -1906
rect 2532 -1940 2566 -1906
rect 2600 -1940 2634 -1906
rect 2668 -1940 2702 -1906
rect 2736 -1940 2770 -1906
rect 2026 -1974 2770 -1940
rect 3026 -1264 3770 -1230
rect 3026 -1298 3060 -1264
rect 3094 -1298 3128 -1264
rect 3162 -1298 3196 -1264
rect 3230 -1298 3264 -1264
rect 3298 -1298 3498 -1264
rect 3532 -1298 3566 -1264
rect 3600 -1298 3634 -1264
rect 3668 -1298 3702 -1264
rect 3736 -1298 3770 -1264
rect 3026 -1331 3770 -1298
rect 3026 -1332 3127 -1331
rect 3026 -1366 3060 -1332
rect 3094 -1366 3127 -1332
rect 3026 -1400 3127 -1366
rect 3669 -1332 3770 -1331
rect 3669 -1366 3702 -1332
rect 3736 -1366 3770 -1332
rect 3026 -1434 3060 -1400
rect 3094 -1434 3127 -1400
rect 3026 -1468 3127 -1434
rect 3026 -1502 3060 -1468
rect 3094 -1502 3127 -1468
rect 3026 -1702 3127 -1502
rect 3026 -1736 3060 -1702
rect 3094 -1736 3127 -1702
rect 3026 -1770 3127 -1736
rect 3026 -1804 3060 -1770
rect 3094 -1804 3127 -1770
rect 3026 -1838 3127 -1804
rect 3189 -1417 3607 -1393
rect 3189 -1451 3213 -1417
rect 3247 -1451 3281 -1417
rect 3315 -1451 3481 -1417
rect 3515 -1451 3549 -1417
rect 3583 -1451 3607 -1417
rect 3189 -1465 3607 -1451
rect 3189 -1485 3261 -1465
rect 3189 -1519 3213 -1485
rect 3247 -1519 3261 -1485
rect 3189 -1685 3261 -1519
rect 3535 -1485 3607 -1465
rect 3535 -1519 3549 -1485
rect 3583 -1519 3607 -1485
rect 3319 -1537 3477 -1523
rect 3319 -1571 3333 -1537
rect 3367 -1551 3429 -1537
rect 3463 -1571 3477 -1537
rect 3319 -1633 3347 -1571
rect 3449 -1633 3477 -1571
rect 3319 -1667 3333 -1633
rect 3367 -1667 3429 -1653
rect 3463 -1667 3477 -1633
rect 3319 -1681 3477 -1667
rect 3189 -1719 3213 -1685
rect 3247 -1719 3261 -1685
rect 3189 -1739 3261 -1719
rect 3535 -1685 3607 -1519
rect 3535 -1719 3549 -1685
rect 3583 -1719 3607 -1685
rect 3535 -1739 3607 -1719
rect 3189 -1753 3607 -1739
rect 3189 -1787 3213 -1753
rect 3247 -1787 3281 -1753
rect 3315 -1787 3481 -1753
rect 3515 -1787 3549 -1753
rect 3583 -1787 3607 -1753
rect 3189 -1811 3607 -1787
rect 3669 -1400 3770 -1366
rect 3669 -1434 3702 -1400
rect 3736 -1434 3770 -1400
rect 3669 -1468 3770 -1434
rect 3669 -1502 3702 -1468
rect 3736 -1502 3770 -1468
rect 3669 -1702 3770 -1502
rect 3669 -1736 3702 -1702
rect 3736 -1736 3770 -1702
rect 3669 -1770 3770 -1736
rect 3669 -1804 3702 -1770
rect 3736 -1804 3770 -1770
rect 3026 -1872 3060 -1838
rect 3094 -1872 3127 -1838
rect 3026 -1873 3127 -1872
rect 3669 -1838 3770 -1804
rect 3669 -1872 3702 -1838
rect 3736 -1872 3770 -1838
rect 3669 -1873 3770 -1872
rect 3026 -1906 3770 -1873
rect 3026 -1940 3060 -1906
rect 3094 -1940 3128 -1906
rect 3162 -1940 3196 -1906
rect 3230 -1940 3264 -1906
rect 3298 -1940 3498 -1906
rect 3532 -1940 3566 -1906
rect 3600 -1940 3634 -1906
rect 3668 -1940 3702 -1906
rect 3736 -1940 3770 -1906
rect 3026 -1974 3770 -1940
rect -974 -2264 -230 -2230
rect -974 -2298 -940 -2264
rect -906 -2298 -872 -2264
rect -838 -2298 -804 -2264
rect -770 -2298 -736 -2264
rect -702 -2298 -502 -2264
rect -468 -2298 -434 -2264
rect -400 -2298 -366 -2264
rect -332 -2298 -298 -2264
rect -264 -2298 -230 -2264
rect -974 -2331 -230 -2298
rect -974 -2332 -873 -2331
rect -974 -2366 -940 -2332
rect -906 -2366 -873 -2332
rect -974 -2400 -873 -2366
rect -331 -2332 -230 -2331
rect -331 -2366 -298 -2332
rect -264 -2366 -230 -2332
rect -974 -2434 -940 -2400
rect -906 -2434 -873 -2400
rect -974 -2468 -873 -2434
rect -974 -2502 -940 -2468
rect -906 -2502 -873 -2468
rect -974 -2702 -873 -2502
rect -974 -2736 -940 -2702
rect -906 -2736 -873 -2702
rect -974 -2770 -873 -2736
rect -974 -2804 -940 -2770
rect -906 -2804 -873 -2770
rect -974 -2838 -873 -2804
rect -811 -2417 -393 -2393
rect -811 -2451 -787 -2417
rect -753 -2451 -719 -2417
rect -685 -2451 -519 -2417
rect -485 -2451 -451 -2417
rect -417 -2451 -393 -2417
rect -811 -2465 -393 -2451
rect -811 -2485 -739 -2465
rect -811 -2519 -787 -2485
rect -753 -2519 -739 -2485
rect -811 -2685 -739 -2519
rect -465 -2485 -393 -2465
rect -465 -2519 -451 -2485
rect -417 -2519 -393 -2485
rect -681 -2537 -523 -2523
rect -681 -2571 -667 -2537
rect -633 -2551 -571 -2537
rect -537 -2571 -523 -2537
rect -681 -2633 -653 -2571
rect -551 -2633 -523 -2571
rect -681 -2667 -667 -2633
rect -633 -2667 -571 -2653
rect -537 -2667 -523 -2633
rect -681 -2681 -523 -2667
rect -811 -2719 -787 -2685
rect -753 -2719 -739 -2685
rect -811 -2739 -739 -2719
rect -465 -2685 -393 -2519
rect -465 -2719 -451 -2685
rect -417 -2719 -393 -2685
rect -465 -2739 -393 -2719
rect -811 -2753 -393 -2739
rect -811 -2787 -787 -2753
rect -753 -2787 -719 -2753
rect -685 -2787 -519 -2753
rect -485 -2787 -451 -2753
rect -417 -2787 -393 -2753
rect -811 -2811 -393 -2787
rect -331 -2400 -230 -2366
rect -331 -2434 -298 -2400
rect -264 -2434 -230 -2400
rect -331 -2468 -230 -2434
rect -331 -2502 -298 -2468
rect -264 -2502 -230 -2468
rect -331 -2702 -230 -2502
rect -331 -2736 -298 -2702
rect -264 -2736 -230 -2702
rect -331 -2770 -230 -2736
rect -331 -2804 -298 -2770
rect -264 -2804 -230 -2770
rect -974 -2872 -940 -2838
rect -906 -2872 -873 -2838
rect -974 -2873 -873 -2872
rect -331 -2838 -230 -2804
rect -331 -2872 -298 -2838
rect -264 -2872 -230 -2838
rect -331 -2873 -230 -2872
rect -974 -2906 -230 -2873
rect -974 -2940 -940 -2906
rect -906 -2940 -872 -2906
rect -838 -2940 -804 -2906
rect -770 -2940 -736 -2906
rect -702 -2940 -502 -2906
rect -468 -2940 -434 -2906
rect -400 -2940 -366 -2906
rect -332 -2940 -298 -2906
rect -264 -2940 -230 -2906
rect -974 -2974 -230 -2940
rect 26 -2264 770 -2230
rect 26 -2298 60 -2264
rect 94 -2298 128 -2264
rect 162 -2298 196 -2264
rect 230 -2298 264 -2264
rect 298 -2298 498 -2264
rect 532 -2298 566 -2264
rect 600 -2298 634 -2264
rect 668 -2298 702 -2264
rect 736 -2298 770 -2264
rect 26 -2331 770 -2298
rect 26 -2332 127 -2331
rect 26 -2366 60 -2332
rect 94 -2366 127 -2332
rect 26 -2400 127 -2366
rect 669 -2332 770 -2331
rect 669 -2366 702 -2332
rect 736 -2366 770 -2332
rect 26 -2434 60 -2400
rect 94 -2434 127 -2400
rect 26 -2468 127 -2434
rect 26 -2502 60 -2468
rect 94 -2502 127 -2468
rect 26 -2702 127 -2502
rect 26 -2736 60 -2702
rect 94 -2736 127 -2702
rect 26 -2770 127 -2736
rect 26 -2804 60 -2770
rect 94 -2804 127 -2770
rect 26 -2838 127 -2804
rect 189 -2417 607 -2393
rect 189 -2451 213 -2417
rect 247 -2451 281 -2417
rect 315 -2451 481 -2417
rect 515 -2451 549 -2417
rect 583 -2451 607 -2417
rect 189 -2465 607 -2451
rect 189 -2485 261 -2465
rect 189 -2519 213 -2485
rect 247 -2519 261 -2485
rect 189 -2685 261 -2519
rect 535 -2485 607 -2465
rect 535 -2519 549 -2485
rect 583 -2519 607 -2485
rect 319 -2537 477 -2523
rect 319 -2571 333 -2537
rect 367 -2551 429 -2537
rect 463 -2571 477 -2537
rect 319 -2633 347 -2571
rect 449 -2633 477 -2571
rect 319 -2667 333 -2633
rect 367 -2667 429 -2653
rect 463 -2667 477 -2633
rect 319 -2681 477 -2667
rect 189 -2719 213 -2685
rect 247 -2719 261 -2685
rect 189 -2739 261 -2719
rect 535 -2685 607 -2519
rect 535 -2719 549 -2685
rect 583 -2719 607 -2685
rect 535 -2739 607 -2719
rect 189 -2753 607 -2739
rect 189 -2787 213 -2753
rect 247 -2787 281 -2753
rect 315 -2787 481 -2753
rect 515 -2787 549 -2753
rect 583 -2787 607 -2753
rect 189 -2811 607 -2787
rect 669 -2400 770 -2366
rect 669 -2434 702 -2400
rect 736 -2434 770 -2400
rect 669 -2468 770 -2434
rect 669 -2502 702 -2468
rect 736 -2502 770 -2468
rect 669 -2702 770 -2502
rect 669 -2736 702 -2702
rect 736 -2736 770 -2702
rect 669 -2770 770 -2736
rect 669 -2804 702 -2770
rect 736 -2804 770 -2770
rect 26 -2872 60 -2838
rect 94 -2872 127 -2838
rect 26 -2873 127 -2872
rect 669 -2838 770 -2804
rect 669 -2872 702 -2838
rect 736 -2872 770 -2838
rect 669 -2873 770 -2872
rect 26 -2906 770 -2873
rect 26 -2940 60 -2906
rect 94 -2940 128 -2906
rect 162 -2940 196 -2906
rect 230 -2940 264 -2906
rect 298 -2940 498 -2906
rect 532 -2940 566 -2906
rect 600 -2940 634 -2906
rect 668 -2940 702 -2906
rect 736 -2940 770 -2906
rect 26 -2974 770 -2940
rect 1026 -2264 1770 -2230
rect 1026 -2298 1060 -2264
rect 1094 -2298 1128 -2264
rect 1162 -2298 1196 -2264
rect 1230 -2298 1264 -2264
rect 1298 -2298 1498 -2264
rect 1532 -2298 1566 -2264
rect 1600 -2298 1634 -2264
rect 1668 -2298 1702 -2264
rect 1736 -2298 1770 -2264
rect 1026 -2331 1770 -2298
rect 1026 -2332 1127 -2331
rect 1026 -2366 1060 -2332
rect 1094 -2366 1127 -2332
rect 1026 -2400 1127 -2366
rect 1669 -2332 1770 -2331
rect 1669 -2366 1702 -2332
rect 1736 -2366 1770 -2332
rect 1026 -2434 1060 -2400
rect 1094 -2434 1127 -2400
rect 1026 -2468 1127 -2434
rect 1026 -2502 1060 -2468
rect 1094 -2502 1127 -2468
rect 1026 -2702 1127 -2502
rect 1026 -2736 1060 -2702
rect 1094 -2736 1127 -2702
rect 1026 -2770 1127 -2736
rect 1026 -2804 1060 -2770
rect 1094 -2804 1127 -2770
rect 1026 -2838 1127 -2804
rect 1189 -2417 1607 -2393
rect 1189 -2451 1213 -2417
rect 1247 -2451 1281 -2417
rect 1315 -2451 1481 -2417
rect 1515 -2451 1549 -2417
rect 1583 -2451 1607 -2417
rect 1189 -2465 1607 -2451
rect 1189 -2485 1261 -2465
rect 1189 -2519 1213 -2485
rect 1247 -2519 1261 -2485
rect 1189 -2685 1261 -2519
rect 1535 -2485 1607 -2465
rect 1535 -2519 1549 -2485
rect 1583 -2519 1607 -2485
rect 1319 -2537 1477 -2523
rect 1319 -2571 1333 -2537
rect 1367 -2551 1429 -2537
rect 1463 -2571 1477 -2537
rect 1319 -2633 1347 -2571
rect 1449 -2633 1477 -2571
rect 1319 -2667 1333 -2633
rect 1367 -2667 1429 -2653
rect 1463 -2667 1477 -2633
rect 1319 -2681 1477 -2667
rect 1189 -2719 1213 -2685
rect 1247 -2719 1261 -2685
rect 1189 -2739 1261 -2719
rect 1535 -2685 1607 -2519
rect 1535 -2719 1549 -2685
rect 1583 -2719 1607 -2685
rect 1535 -2739 1607 -2719
rect 1189 -2753 1607 -2739
rect 1189 -2787 1213 -2753
rect 1247 -2787 1281 -2753
rect 1315 -2787 1481 -2753
rect 1515 -2787 1549 -2753
rect 1583 -2787 1607 -2753
rect 1189 -2811 1607 -2787
rect 1669 -2400 1770 -2366
rect 1669 -2434 1702 -2400
rect 1736 -2434 1770 -2400
rect 1669 -2468 1770 -2434
rect 1669 -2502 1702 -2468
rect 1736 -2502 1770 -2468
rect 1669 -2702 1770 -2502
rect 1669 -2736 1702 -2702
rect 1736 -2736 1770 -2702
rect 1669 -2770 1770 -2736
rect 1669 -2804 1702 -2770
rect 1736 -2804 1770 -2770
rect 1026 -2872 1060 -2838
rect 1094 -2872 1127 -2838
rect 1026 -2873 1127 -2872
rect 1669 -2838 1770 -2804
rect 1669 -2872 1702 -2838
rect 1736 -2872 1770 -2838
rect 1669 -2873 1770 -2872
rect 1026 -2906 1770 -2873
rect 1026 -2940 1060 -2906
rect 1094 -2940 1128 -2906
rect 1162 -2940 1196 -2906
rect 1230 -2940 1264 -2906
rect 1298 -2940 1498 -2906
rect 1532 -2940 1566 -2906
rect 1600 -2940 1634 -2906
rect 1668 -2940 1702 -2906
rect 1736 -2940 1770 -2906
rect 1026 -2974 1770 -2940
rect 2026 -2264 2770 -2230
rect 2026 -2298 2060 -2264
rect 2094 -2298 2128 -2264
rect 2162 -2298 2196 -2264
rect 2230 -2298 2264 -2264
rect 2298 -2298 2498 -2264
rect 2532 -2298 2566 -2264
rect 2600 -2298 2634 -2264
rect 2668 -2298 2702 -2264
rect 2736 -2298 2770 -2264
rect 2026 -2331 2770 -2298
rect 2026 -2332 2127 -2331
rect 2026 -2366 2060 -2332
rect 2094 -2366 2127 -2332
rect 2026 -2400 2127 -2366
rect 2669 -2332 2770 -2331
rect 2669 -2366 2702 -2332
rect 2736 -2366 2770 -2332
rect 2026 -2434 2060 -2400
rect 2094 -2434 2127 -2400
rect 2026 -2468 2127 -2434
rect 2026 -2502 2060 -2468
rect 2094 -2502 2127 -2468
rect 2026 -2702 2127 -2502
rect 2026 -2736 2060 -2702
rect 2094 -2736 2127 -2702
rect 2026 -2770 2127 -2736
rect 2026 -2804 2060 -2770
rect 2094 -2804 2127 -2770
rect 2026 -2838 2127 -2804
rect 2189 -2417 2607 -2393
rect 2189 -2451 2213 -2417
rect 2247 -2451 2281 -2417
rect 2315 -2451 2481 -2417
rect 2515 -2451 2549 -2417
rect 2583 -2451 2607 -2417
rect 2189 -2465 2607 -2451
rect 2189 -2485 2261 -2465
rect 2189 -2519 2213 -2485
rect 2247 -2519 2261 -2485
rect 2189 -2685 2261 -2519
rect 2535 -2485 2607 -2465
rect 2535 -2519 2549 -2485
rect 2583 -2519 2607 -2485
rect 2319 -2537 2477 -2523
rect 2319 -2571 2333 -2537
rect 2367 -2551 2429 -2537
rect 2463 -2571 2477 -2537
rect 2319 -2633 2347 -2571
rect 2449 -2633 2477 -2571
rect 2319 -2667 2333 -2633
rect 2367 -2667 2429 -2653
rect 2463 -2667 2477 -2633
rect 2319 -2681 2477 -2667
rect 2189 -2719 2213 -2685
rect 2247 -2719 2261 -2685
rect 2189 -2739 2261 -2719
rect 2535 -2685 2607 -2519
rect 2535 -2719 2549 -2685
rect 2583 -2719 2607 -2685
rect 2535 -2739 2607 -2719
rect 2189 -2753 2607 -2739
rect 2189 -2787 2213 -2753
rect 2247 -2787 2281 -2753
rect 2315 -2787 2481 -2753
rect 2515 -2787 2549 -2753
rect 2583 -2787 2607 -2753
rect 2189 -2811 2607 -2787
rect 2669 -2400 2770 -2366
rect 2669 -2434 2702 -2400
rect 2736 -2434 2770 -2400
rect 2669 -2468 2770 -2434
rect 2669 -2502 2702 -2468
rect 2736 -2502 2770 -2468
rect 2669 -2702 2770 -2502
rect 2669 -2736 2702 -2702
rect 2736 -2736 2770 -2702
rect 2669 -2770 2770 -2736
rect 2669 -2804 2702 -2770
rect 2736 -2804 2770 -2770
rect 2026 -2872 2060 -2838
rect 2094 -2872 2127 -2838
rect 2026 -2873 2127 -2872
rect 2669 -2838 2770 -2804
rect 2669 -2872 2702 -2838
rect 2736 -2872 2770 -2838
rect 2669 -2873 2770 -2872
rect 2026 -2906 2770 -2873
rect 2026 -2940 2060 -2906
rect 2094 -2940 2128 -2906
rect 2162 -2940 2196 -2906
rect 2230 -2940 2264 -2906
rect 2298 -2940 2498 -2906
rect 2532 -2940 2566 -2906
rect 2600 -2940 2634 -2906
rect 2668 -2940 2702 -2906
rect 2736 -2940 2770 -2906
rect 2026 -2974 2770 -2940
rect 3026 -2264 3770 -2230
rect 3026 -2298 3060 -2264
rect 3094 -2298 3128 -2264
rect 3162 -2298 3196 -2264
rect 3230 -2298 3264 -2264
rect 3298 -2298 3498 -2264
rect 3532 -2298 3566 -2264
rect 3600 -2298 3634 -2264
rect 3668 -2298 3702 -2264
rect 3736 -2298 3770 -2264
rect 3026 -2331 3770 -2298
rect 3026 -2332 3127 -2331
rect 3026 -2366 3060 -2332
rect 3094 -2366 3127 -2332
rect 3026 -2400 3127 -2366
rect 3669 -2332 3770 -2331
rect 3669 -2366 3702 -2332
rect 3736 -2366 3770 -2332
rect 3026 -2434 3060 -2400
rect 3094 -2434 3127 -2400
rect 3026 -2468 3127 -2434
rect 3026 -2502 3060 -2468
rect 3094 -2502 3127 -2468
rect 3026 -2702 3127 -2502
rect 3026 -2736 3060 -2702
rect 3094 -2736 3127 -2702
rect 3026 -2770 3127 -2736
rect 3026 -2804 3060 -2770
rect 3094 -2804 3127 -2770
rect 3026 -2838 3127 -2804
rect 3189 -2417 3607 -2393
rect 3189 -2451 3213 -2417
rect 3247 -2451 3281 -2417
rect 3315 -2451 3481 -2417
rect 3515 -2451 3549 -2417
rect 3583 -2451 3607 -2417
rect 3189 -2465 3607 -2451
rect 3189 -2485 3261 -2465
rect 3189 -2519 3213 -2485
rect 3247 -2519 3261 -2485
rect 3189 -2685 3261 -2519
rect 3535 -2485 3607 -2465
rect 3535 -2519 3549 -2485
rect 3583 -2519 3607 -2485
rect 3319 -2537 3477 -2523
rect 3319 -2571 3333 -2537
rect 3367 -2551 3429 -2537
rect 3463 -2571 3477 -2537
rect 3319 -2633 3347 -2571
rect 3449 -2633 3477 -2571
rect 3319 -2667 3333 -2633
rect 3367 -2667 3429 -2653
rect 3463 -2667 3477 -2633
rect 3319 -2681 3477 -2667
rect 3189 -2719 3213 -2685
rect 3247 -2719 3261 -2685
rect 3189 -2739 3261 -2719
rect 3535 -2685 3607 -2519
rect 3535 -2719 3549 -2685
rect 3583 -2719 3607 -2685
rect 3535 -2739 3607 -2719
rect 3189 -2753 3607 -2739
rect 3189 -2787 3213 -2753
rect 3247 -2787 3281 -2753
rect 3315 -2787 3481 -2753
rect 3515 -2787 3549 -2753
rect 3583 -2787 3607 -2753
rect 3189 -2811 3607 -2787
rect 3669 -2400 3770 -2366
rect 3669 -2434 3702 -2400
rect 3736 -2434 3770 -2400
rect 3669 -2468 3770 -2434
rect 3669 -2502 3702 -2468
rect 3736 -2502 3770 -2468
rect 3669 -2702 3770 -2502
rect 3669 -2736 3702 -2702
rect 3736 -2736 3770 -2702
rect 3669 -2770 3770 -2736
rect 3669 -2804 3702 -2770
rect 3736 -2804 3770 -2770
rect 3026 -2872 3060 -2838
rect 3094 -2872 3127 -2838
rect 3026 -2873 3127 -2872
rect 3669 -2838 3770 -2804
rect 3669 -2872 3702 -2838
rect 3736 -2872 3770 -2838
rect 3669 -2873 3770 -2872
rect 3026 -2906 3770 -2873
rect 3026 -2940 3060 -2906
rect 3094 -2940 3128 -2906
rect 3162 -2940 3196 -2906
rect 3230 -2940 3264 -2906
rect 3298 -2940 3498 -2906
rect 3532 -2940 3566 -2906
rect 3600 -2940 3634 -2906
rect 3668 -2940 3702 -2906
rect 3736 -2940 3770 -2906
rect 3026 -2974 3770 -2940
<< viali >>
rect -3667 1449 -3633 1463
rect -3571 1449 -3537 1463
rect -3667 1429 -3653 1449
rect -3653 1429 -3633 1449
rect -3571 1429 -3551 1449
rect -3551 1429 -3537 1449
rect -3667 1347 -3653 1367
rect -3653 1347 -3633 1367
rect -3571 1347 -3551 1367
rect -3551 1347 -3537 1367
rect -3667 1333 -3633 1347
rect -3571 1333 -3537 1347
rect -2667 1449 -2633 1463
rect -2571 1449 -2537 1463
rect -2667 1429 -2653 1449
rect -2653 1429 -2633 1449
rect -2571 1429 -2551 1449
rect -2551 1429 -2537 1449
rect -2667 1347 -2653 1367
rect -2653 1347 -2633 1367
rect -2571 1347 -2551 1367
rect -2551 1347 -2537 1367
rect -2667 1333 -2633 1347
rect -2571 1333 -2537 1347
rect -1667 1449 -1633 1463
rect -1571 1449 -1537 1463
rect -1667 1429 -1653 1449
rect -1653 1429 -1633 1449
rect -1571 1429 -1551 1449
rect -1551 1429 -1537 1449
rect -1667 1347 -1653 1367
rect -1653 1347 -1633 1367
rect -1571 1347 -1551 1367
rect -1551 1347 -1537 1367
rect -1667 1333 -1633 1347
rect -1571 1333 -1537 1347
rect -667 1449 -633 1463
rect -571 1449 -537 1463
rect -667 1429 -653 1449
rect -653 1429 -633 1449
rect -571 1429 -551 1449
rect -551 1429 -537 1449
rect -667 1347 -653 1367
rect -653 1347 -633 1367
rect -571 1347 -551 1367
rect -551 1347 -537 1367
rect -667 1333 -633 1347
rect -571 1333 -537 1347
rect 333 1449 367 1463
rect 429 1449 463 1463
rect 333 1429 347 1449
rect 347 1429 367 1449
rect 429 1429 449 1449
rect 449 1429 463 1449
rect 333 1347 347 1367
rect 347 1347 367 1367
rect 429 1347 449 1367
rect 449 1347 463 1367
rect 333 1333 367 1347
rect 429 1333 463 1347
rect 1333 1449 1367 1463
rect 1429 1449 1463 1463
rect 1333 1429 1347 1449
rect 1347 1429 1367 1449
rect 1429 1429 1449 1449
rect 1449 1429 1463 1449
rect 1333 1347 1347 1367
rect 1347 1347 1367 1367
rect 1429 1347 1449 1367
rect 1449 1347 1463 1367
rect 1333 1333 1367 1347
rect 1429 1333 1463 1347
rect 2333 1449 2367 1463
rect 2429 1449 2463 1463
rect 2333 1429 2347 1449
rect 2347 1429 2367 1449
rect 2429 1429 2449 1449
rect 2449 1429 2463 1449
rect 2333 1347 2347 1367
rect 2347 1347 2367 1367
rect 2429 1347 2449 1367
rect 2449 1347 2463 1367
rect 2333 1333 2367 1347
rect 2429 1333 2463 1347
rect 3333 1449 3367 1463
rect 3429 1449 3463 1463
rect 3333 1429 3347 1449
rect 3347 1429 3367 1449
rect 3429 1429 3449 1449
rect 3449 1429 3463 1449
rect 3333 1347 3347 1367
rect 3347 1347 3367 1367
rect 3429 1347 3449 1367
rect 3449 1347 3463 1367
rect 3333 1333 3367 1347
rect 3429 1333 3463 1347
rect -3667 449 -3633 463
rect -3571 449 -3537 463
rect -3667 429 -3653 449
rect -3653 429 -3633 449
rect -3571 429 -3551 449
rect -3551 429 -3537 449
rect -3667 347 -3653 367
rect -3653 347 -3633 367
rect -3571 347 -3551 367
rect -3551 347 -3537 367
rect -3667 333 -3633 347
rect -3571 333 -3537 347
rect -2667 449 -2633 463
rect -2571 449 -2537 463
rect -2667 429 -2653 449
rect -2653 429 -2633 449
rect -2571 429 -2551 449
rect -2551 429 -2537 449
rect -2667 347 -2653 367
rect -2653 347 -2633 367
rect -2571 347 -2551 367
rect -2551 347 -2537 367
rect -2667 333 -2633 347
rect -2571 333 -2537 347
rect -1667 449 -1633 463
rect -1571 449 -1537 463
rect -1667 429 -1653 449
rect -1653 429 -1633 449
rect -1571 429 -1551 449
rect -1551 429 -1537 449
rect -1667 347 -1653 367
rect -1653 347 -1633 367
rect -1571 347 -1551 367
rect -1551 347 -1537 367
rect -1667 333 -1633 347
rect -1571 333 -1537 347
rect -667 449 -633 463
rect -571 449 -537 463
rect -667 429 -653 449
rect -653 429 -633 449
rect -571 429 -551 449
rect -551 429 -537 449
rect -667 347 -653 367
rect -653 347 -633 367
rect -571 347 -551 367
rect -551 347 -537 367
rect -667 333 -633 347
rect -571 333 -537 347
rect 1333 449 1367 463
rect 1429 449 1463 463
rect 1333 429 1347 449
rect 1347 429 1367 449
rect 1429 429 1449 449
rect 1449 429 1463 449
rect 1333 347 1347 367
rect 1347 347 1367 367
rect 1429 347 1449 367
rect 1449 347 1463 367
rect 1333 333 1367 347
rect 1429 333 1463 347
rect 2333 449 2367 463
rect 2429 449 2463 463
rect 2333 429 2347 449
rect 2347 429 2367 449
rect 2429 429 2449 449
rect 2449 429 2463 449
rect 2333 347 2347 367
rect 2347 347 2367 367
rect 2429 347 2449 367
rect 2449 347 2463 367
rect 2333 333 2367 347
rect 2429 333 2463 347
rect 3333 449 3367 463
rect 3429 449 3463 463
rect 3333 429 3347 449
rect 3347 429 3367 449
rect 3429 429 3449 449
rect 3449 429 3463 449
rect 3333 347 3347 367
rect 3347 347 3367 367
rect 3429 347 3449 367
rect 3449 347 3463 367
rect 3333 333 3367 347
rect 3429 333 3463 347
rect -3667 -551 -3633 -537
rect -3571 -551 -3537 -537
rect -3667 -571 -3653 -551
rect -3653 -571 -3633 -551
rect -3571 -571 -3551 -551
rect -3551 -571 -3537 -551
rect -3667 -653 -3653 -633
rect -3653 -653 -3633 -633
rect -3571 -653 -3551 -633
rect -3551 -653 -3537 -633
rect -3667 -667 -3633 -653
rect -3571 -667 -3537 -653
rect -2667 -551 -2633 -537
rect -2571 -551 -2537 -537
rect -2667 -571 -2653 -551
rect -2653 -571 -2633 -551
rect -2571 -571 -2551 -551
rect -2551 -571 -2537 -551
rect -2667 -653 -2653 -633
rect -2653 -653 -2633 -633
rect -2571 -653 -2551 -633
rect -2551 -653 -2537 -633
rect -2667 -667 -2633 -653
rect -2571 -667 -2537 -653
rect -1667 -551 -1633 -537
rect -1571 -551 -1537 -537
rect -1667 -571 -1653 -551
rect -1653 -571 -1633 -551
rect -1571 -571 -1551 -551
rect -1551 -571 -1537 -551
rect -1667 -653 -1653 -633
rect -1653 -653 -1633 -633
rect -1571 -653 -1551 -633
rect -1551 -653 -1537 -633
rect -1667 -667 -1633 -653
rect -1571 -667 -1537 -653
rect -667 -551 -633 -537
rect -571 -551 -537 -537
rect -667 -571 -653 -551
rect -653 -571 -633 -551
rect -571 -571 -551 -551
rect -551 -571 -537 -551
rect -667 -653 -653 -633
rect -653 -653 -633 -633
rect -571 -653 -551 -633
rect -551 -653 -537 -633
rect -667 -667 -633 -653
rect -571 -667 -537 -653
rect 333 -551 367 -537
rect 429 -551 463 -537
rect 333 -571 347 -551
rect 347 -571 367 -551
rect 429 -571 449 -551
rect 449 -571 463 -551
rect 333 -653 347 -633
rect 347 -653 367 -633
rect 429 -653 449 -633
rect 449 -653 463 -633
rect 333 -667 367 -653
rect 429 -667 463 -653
rect 1333 -551 1367 -537
rect 1429 -551 1463 -537
rect 1333 -571 1347 -551
rect 1347 -571 1367 -551
rect 1429 -571 1449 -551
rect 1449 -571 1463 -551
rect 1333 -653 1347 -633
rect 1347 -653 1367 -633
rect 1429 -653 1449 -633
rect 1449 -653 1463 -633
rect 1333 -667 1367 -653
rect 1429 -667 1463 -653
rect 2333 -551 2367 -537
rect 2429 -551 2463 -537
rect 2333 -571 2347 -551
rect 2347 -571 2367 -551
rect 2429 -571 2449 -551
rect 2449 -571 2463 -551
rect 2333 -653 2347 -633
rect 2347 -653 2367 -633
rect 2429 -653 2449 -633
rect 2449 -653 2463 -633
rect 2333 -667 2367 -653
rect 2429 -667 2463 -653
rect 3333 -551 3367 -537
rect 3429 -551 3463 -537
rect 3333 -571 3347 -551
rect 3347 -571 3367 -551
rect 3429 -571 3449 -551
rect 3449 -571 3463 -551
rect 3333 -653 3347 -633
rect 3347 -653 3367 -633
rect 3429 -653 3449 -633
rect 3449 -653 3463 -633
rect 3333 -667 3367 -653
rect 3429 -667 3463 -653
rect -667 -1551 -633 -1537
rect -571 -1551 -537 -1537
rect -667 -1571 -653 -1551
rect -653 -1571 -633 -1551
rect -571 -1571 -551 -1551
rect -551 -1571 -537 -1551
rect -667 -1653 -653 -1633
rect -653 -1653 -633 -1633
rect -571 -1653 -551 -1633
rect -551 -1653 -537 -1633
rect -667 -1667 -633 -1653
rect -571 -1667 -537 -1653
rect 333 -1551 367 -1537
rect 429 -1551 463 -1537
rect 333 -1571 347 -1551
rect 347 -1571 367 -1551
rect 429 -1571 449 -1551
rect 449 -1571 463 -1551
rect 333 -1653 347 -1633
rect 347 -1653 367 -1633
rect 429 -1653 449 -1633
rect 449 -1653 463 -1633
rect 333 -1667 367 -1653
rect 429 -1667 463 -1653
rect 1333 -1551 1367 -1537
rect 1429 -1551 1463 -1537
rect 1333 -1571 1347 -1551
rect 1347 -1571 1367 -1551
rect 1429 -1571 1449 -1551
rect 1449 -1571 1463 -1551
rect 1333 -1653 1347 -1633
rect 1347 -1653 1367 -1633
rect 1429 -1653 1449 -1633
rect 1449 -1653 1463 -1633
rect 1333 -1667 1367 -1653
rect 1429 -1667 1463 -1653
rect 2333 -1551 2367 -1537
rect 2429 -1551 2463 -1537
rect 2333 -1571 2347 -1551
rect 2347 -1571 2367 -1551
rect 2429 -1571 2449 -1551
rect 2449 -1571 2463 -1551
rect 2333 -1653 2347 -1633
rect 2347 -1653 2367 -1633
rect 2429 -1653 2449 -1633
rect 2449 -1653 2463 -1633
rect 2333 -1667 2367 -1653
rect 2429 -1667 2463 -1653
rect 3333 -1551 3367 -1537
rect 3429 -1551 3463 -1537
rect 3333 -1571 3347 -1551
rect 3347 -1571 3367 -1551
rect 3429 -1571 3449 -1551
rect 3449 -1571 3463 -1551
rect 3333 -1653 3347 -1633
rect 3347 -1653 3367 -1633
rect 3429 -1653 3449 -1633
rect 3449 -1653 3463 -1633
rect 3333 -1667 3367 -1653
rect 3429 -1667 3463 -1653
rect -667 -2551 -633 -2537
rect -571 -2551 -537 -2537
rect -667 -2571 -653 -2551
rect -653 -2571 -633 -2551
rect -571 -2571 -551 -2551
rect -551 -2571 -537 -2551
rect -667 -2653 -653 -2633
rect -653 -2653 -633 -2633
rect -571 -2653 -551 -2633
rect -551 -2653 -537 -2633
rect -667 -2667 -633 -2653
rect -571 -2667 -537 -2653
rect 333 -2551 367 -2537
rect 429 -2551 463 -2537
rect 333 -2571 347 -2551
rect 347 -2571 367 -2551
rect 429 -2571 449 -2551
rect 449 -2571 463 -2551
rect 333 -2653 347 -2633
rect 347 -2653 367 -2633
rect 429 -2653 449 -2633
rect 449 -2653 463 -2633
rect 333 -2667 367 -2653
rect 429 -2667 463 -2653
rect 1333 -2551 1367 -2537
rect 1429 -2551 1463 -2537
rect 1333 -2571 1347 -2551
rect 1347 -2571 1367 -2551
rect 1429 -2571 1449 -2551
rect 1449 -2571 1463 -2551
rect 1333 -2653 1347 -2633
rect 1347 -2653 1367 -2633
rect 1429 -2653 1449 -2633
rect 1449 -2653 1463 -2633
rect 1333 -2667 1367 -2653
rect 1429 -2667 1463 -2653
rect 2333 -2551 2367 -2537
rect 2429 -2551 2463 -2537
rect 2333 -2571 2347 -2551
rect 2347 -2571 2367 -2551
rect 2429 -2571 2449 -2551
rect 2449 -2571 2463 -2551
rect 2333 -2653 2347 -2633
rect 2347 -2653 2367 -2633
rect 2429 -2653 2449 -2633
rect 2449 -2653 2463 -2633
rect 2333 -2667 2367 -2653
rect 2429 -2667 2463 -2653
rect 3333 -2551 3367 -2537
rect 3429 -2551 3463 -2537
rect 3333 -2571 3347 -2551
rect 3347 -2571 3367 -2551
rect 3429 -2571 3449 -2551
rect 3449 -2571 3463 -2551
rect 3333 -2653 3347 -2633
rect 3347 -2653 3367 -2633
rect 3429 -2653 3449 -2633
rect 3449 -2653 3463 -2633
rect 3333 -2667 3367 -2653
rect 3429 -2667 3463 -2653
<< metal1 >>
rect -3685 1463 -3519 1481
rect -3685 1429 -3667 1463
rect -3633 1429 -3571 1463
rect -3537 1429 -3519 1463
rect -3685 1367 -3519 1429
rect -3685 1333 -3667 1367
rect -3633 1333 -3571 1367
rect -3537 1333 -3519 1367
rect -3685 1315 -3519 1333
rect -2685 1463 -2519 1481
rect -2685 1429 -2667 1463
rect -2633 1429 -2571 1463
rect -2537 1429 -2519 1463
rect -2685 1367 -2519 1429
rect -2685 1333 -2667 1367
rect -2633 1333 -2571 1367
rect -2537 1333 -2519 1367
rect -2685 1315 -2519 1333
rect -1685 1463 -1519 1481
rect -1685 1429 -1667 1463
rect -1633 1429 -1571 1463
rect -1537 1429 -1519 1463
rect -1685 1367 -1519 1429
rect -1685 1333 -1667 1367
rect -1633 1333 -1571 1367
rect -1537 1333 -1519 1367
rect -1685 1315 -1519 1333
rect -685 1463 -519 1481
rect -685 1429 -667 1463
rect -633 1429 -571 1463
rect -537 1429 -519 1463
rect -685 1367 -519 1429
rect -685 1333 -667 1367
rect -633 1333 -571 1367
rect -537 1333 -519 1367
rect -685 1315 -519 1333
rect 315 1463 481 1481
rect 315 1429 333 1463
rect 367 1429 429 1463
rect 463 1429 481 1463
rect 315 1367 481 1429
rect 315 1333 333 1367
rect 367 1333 429 1367
rect 463 1333 481 1367
rect 315 1315 481 1333
rect 1315 1463 1481 1481
rect 1315 1429 1333 1463
rect 1367 1429 1429 1463
rect 1463 1429 1481 1463
rect 1315 1367 1481 1429
rect 1315 1333 1333 1367
rect 1367 1333 1429 1367
rect 1463 1333 1481 1367
rect 1315 1315 1481 1333
rect 2315 1463 2481 1481
rect 2315 1429 2333 1463
rect 2367 1429 2429 1463
rect 2463 1429 2481 1463
rect 2315 1367 2481 1429
rect 2315 1333 2333 1367
rect 2367 1333 2429 1367
rect 2463 1333 2481 1367
rect 2315 1315 2481 1333
rect 3315 1463 3481 1481
rect 3315 1429 3333 1463
rect 3367 1429 3429 1463
rect 3463 1429 3481 1463
rect 3315 1367 3481 1429
rect 3315 1333 3333 1367
rect 3367 1333 3429 1367
rect 3463 1333 3481 1367
rect 3315 1315 3481 1333
rect -3685 463 -3519 481
rect -3685 429 -3667 463
rect -3633 429 -3571 463
rect -3537 429 -3519 463
rect -3685 367 -3519 429
rect -3685 333 -3667 367
rect -3633 333 -3571 367
rect -3537 333 -3519 367
rect -3685 315 -3519 333
rect -2685 463 -2519 481
rect -2685 429 -2667 463
rect -2633 429 -2571 463
rect -2537 429 -2519 463
rect -2685 367 -2519 429
rect -2685 333 -2667 367
rect -2633 333 -2571 367
rect -2537 333 -2519 367
rect -2685 315 -2519 333
rect -1685 463 -1519 481
rect -1685 429 -1667 463
rect -1633 429 -1571 463
rect -1537 429 -1519 463
rect -1685 367 -1519 429
rect -1685 333 -1667 367
rect -1633 333 -1571 367
rect -1537 333 -1519 367
rect -1685 315 -1519 333
rect -685 463 -519 481
rect -685 429 -667 463
rect -633 429 -571 463
rect -537 429 -519 463
rect -685 367 -519 429
rect -685 333 -667 367
rect -633 333 -571 367
rect -537 333 -519 367
rect -685 315 -519 333
rect 1315 463 1481 481
rect 1315 429 1333 463
rect 1367 429 1429 463
rect 1463 429 1481 463
rect 1315 367 1481 429
rect 1315 333 1333 367
rect 1367 333 1429 367
rect 1463 333 1481 367
rect 1315 315 1481 333
rect 2315 463 2481 481
rect 2315 429 2333 463
rect 2367 429 2429 463
rect 2463 429 2481 463
rect 2315 367 2481 429
rect 2315 333 2333 367
rect 2367 333 2429 367
rect 2463 333 2481 367
rect 2315 315 2481 333
rect 3315 463 3481 481
rect 3315 429 3333 463
rect 3367 429 3429 463
rect 3463 429 3481 463
rect 3315 367 3481 429
rect 3315 333 3333 367
rect 3367 333 3429 367
rect 3463 333 3481 367
rect 3315 315 3481 333
rect -3685 -537 -3519 -519
rect -3685 -571 -3667 -537
rect -3633 -571 -3571 -537
rect -3537 -571 -3519 -537
rect -3685 -633 -3519 -571
rect -3685 -667 -3667 -633
rect -3633 -667 -3571 -633
rect -3537 -667 -3519 -633
rect -3685 -685 -3519 -667
rect -2685 -537 -2519 -519
rect -2685 -571 -2667 -537
rect -2633 -571 -2571 -537
rect -2537 -571 -2519 -537
rect -2685 -633 -2519 -571
rect -2685 -667 -2667 -633
rect -2633 -667 -2571 -633
rect -2537 -667 -2519 -633
rect -2685 -685 -2519 -667
rect -1685 -537 -1519 -519
rect -1685 -571 -1667 -537
rect -1633 -571 -1571 -537
rect -1537 -571 -1519 -537
rect -1685 -633 -1519 -571
rect -1685 -667 -1667 -633
rect -1633 -667 -1571 -633
rect -1537 -667 -1519 -633
rect -1685 -685 -1519 -667
rect -685 -537 -519 -519
rect -685 -571 -667 -537
rect -633 -571 -571 -537
rect -537 -571 -519 -537
rect -685 -633 -519 -571
rect -685 -667 -667 -633
rect -633 -667 -571 -633
rect -537 -667 -519 -633
rect -685 -685 -519 -667
rect 315 -537 481 -519
rect 315 -571 333 -537
rect 367 -571 429 -537
rect 463 -571 481 -537
rect 315 -633 481 -571
rect 315 -667 333 -633
rect 367 -667 429 -633
rect 463 -667 481 -633
rect 315 -685 481 -667
rect 1315 -537 1481 -519
rect 1315 -571 1333 -537
rect 1367 -571 1429 -537
rect 1463 -571 1481 -537
rect 1315 -633 1481 -571
rect 1315 -667 1333 -633
rect 1367 -667 1429 -633
rect 1463 -667 1481 -633
rect 1315 -685 1481 -667
rect 2315 -537 2481 -519
rect 2315 -571 2333 -537
rect 2367 -571 2429 -537
rect 2463 -571 2481 -537
rect 2315 -633 2481 -571
rect 2315 -667 2333 -633
rect 2367 -667 2429 -633
rect 2463 -667 2481 -633
rect 2315 -685 2481 -667
rect 3315 -537 3481 -519
rect 3315 -571 3333 -537
rect 3367 -571 3429 -537
rect 3463 -571 3481 -537
rect 3315 -633 3481 -571
rect 3315 -667 3333 -633
rect 3367 -667 3429 -633
rect 3463 -667 3481 -633
rect 3315 -685 3481 -667
rect -685 -1537 -519 -1519
rect -685 -1571 -667 -1537
rect -633 -1571 -571 -1537
rect -537 -1571 -519 -1537
rect -685 -1633 -519 -1571
rect -685 -1667 -667 -1633
rect -633 -1667 -571 -1633
rect -537 -1667 -519 -1633
rect -685 -1685 -519 -1667
rect 315 -1537 481 -1519
rect 315 -1571 333 -1537
rect 367 -1571 429 -1537
rect 463 -1571 481 -1537
rect 315 -1633 481 -1571
rect 315 -1667 333 -1633
rect 367 -1667 429 -1633
rect 463 -1667 481 -1633
rect 315 -1685 481 -1667
rect 1315 -1537 1481 -1519
rect 1315 -1571 1333 -1537
rect 1367 -1571 1429 -1537
rect 1463 -1571 1481 -1537
rect 1315 -1633 1481 -1571
rect 1315 -1667 1333 -1633
rect 1367 -1667 1429 -1633
rect 1463 -1667 1481 -1633
rect 1315 -1685 1481 -1667
rect 2315 -1537 2481 -1519
rect 2315 -1571 2333 -1537
rect 2367 -1571 2429 -1537
rect 2463 -1571 2481 -1537
rect 2315 -1633 2481 -1571
rect 2315 -1667 2333 -1633
rect 2367 -1667 2429 -1633
rect 2463 -1667 2481 -1633
rect 2315 -1685 2481 -1667
rect 3315 -1537 3481 -1519
rect 3315 -1571 3333 -1537
rect 3367 -1571 3429 -1537
rect 3463 -1571 3481 -1537
rect 3315 -1633 3481 -1571
rect 3315 -1667 3333 -1633
rect 3367 -1667 3429 -1633
rect 3463 -1667 3481 -1633
rect 3315 -1685 3481 -1667
rect -685 -2537 -519 -2519
rect -685 -2571 -667 -2537
rect -633 -2571 -571 -2537
rect -537 -2571 -519 -2537
rect -685 -2633 -519 -2571
rect -685 -2667 -667 -2633
rect -633 -2667 -571 -2633
rect -537 -2667 -519 -2633
rect -685 -2685 -519 -2667
rect 315 -2537 481 -2519
rect 315 -2571 333 -2537
rect 367 -2571 429 -2537
rect 463 -2571 481 -2537
rect 315 -2633 481 -2571
rect 315 -2667 333 -2633
rect 367 -2667 429 -2633
rect 463 -2667 481 -2633
rect 315 -2685 481 -2667
rect 1315 -2537 1481 -2519
rect 1315 -2571 1333 -2537
rect 1367 -2571 1429 -2537
rect 1463 -2571 1481 -2537
rect 1315 -2633 1481 -2571
rect 1315 -2667 1333 -2633
rect 1367 -2667 1429 -2633
rect 1463 -2667 1481 -2633
rect 1315 -2685 1481 -2667
rect 2315 -2537 2481 -2519
rect 2315 -2571 2333 -2537
rect 2367 -2571 2429 -2537
rect 2463 -2571 2481 -2537
rect 2315 -2633 2481 -2571
rect 2315 -2667 2333 -2633
rect 2367 -2667 2429 -2633
rect 2463 -2667 2481 -2633
rect 2315 -2685 2481 -2667
rect 3315 -2537 3481 -2519
rect 3315 -2571 3333 -2537
rect 3367 -2571 3429 -2537
rect 3463 -2571 3481 -2537
rect 3315 -2633 3481 -2571
rect 3315 -2667 3333 -2633
rect 3367 -2667 3429 -2633
rect 3463 -2667 3481 -2633
rect 3315 -2685 3481 -2667
<< comment >>
rect -3974 1783 -3973 1796
tri -3973 1783 -3969 1787 se
tri -3235 1783 -3231 1787 sw
rect -3231 1783 -3230 1796
rect -3974 1782 -3629 1783
rect -3576 1782 -3230 1783
rect -3974 1770 -3973 1782
tri -3973 1778 -3969 1782 ne
tri -3235 1778 -3231 1782 nw
rect -3231 1770 -3230 1782
rect -2974 1783 -2973 1796
tri -2973 1783 -2969 1787 se
tri -2235 1783 -2231 1787 sw
rect -2231 1783 -2230 1796
rect -2974 1782 -2629 1783
rect -2576 1782 -2230 1783
rect -2974 1770 -2973 1782
tri -2973 1778 -2969 1782 ne
tri -2235 1778 -2231 1782 nw
rect -2231 1770 -2230 1782
rect -1974 1783 -1973 1796
tri -1973 1783 -1969 1787 se
tri -1235 1783 -1231 1787 sw
rect -1231 1783 -1230 1796
rect -1974 1782 -1629 1783
rect -1576 1782 -1230 1783
rect -1974 1770 -1973 1782
tri -1973 1778 -1969 1782 ne
tri -1235 1778 -1231 1782 nw
rect -1231 1770 -1230 1782
rect -974 1783 -973 1796
tri -973 1783 -969 1787 se
tri -235 1783 -231 1787 sw
rect -231 1783 -230 1796
rect -974 1782 -629 1783
rect -576 1782 -230 1783
rect -974 1770 -973 1782
tri -973 1778 -969 1782 ne
tri -235 1778 -231 1782 nw
rect -231 1770 -230 1782
rect 26 1783 27 1796
tri 27 1783 31 1787 se
tri 765 1783 769 1787 sw
rect 769 1783 770 1796
rect 26 1782 371 1783
rect 424 1782 770 1783
rect 26 1770 27 1782
tri 27 1778 31 1782 ne
tri 765 1778 769 1782 nw
rect 769 1770 770 1782
rect 1026 1783 1027 1796
tri 1027 1783 1031 1787 se
tri 1765 1783 1769 1787 sw
rect 1769 1783 1770 1796
rect 1026 1782 1371 1783
rect 1424 1782 1770 1783
rect 1026 1770 1027 1782
tri 1027 1778 1031 1782 ne
tri 1765 1778 1769 1782 nw
rect 1769 1770 1770 1782
rect 2026 1783 2027 1796
tri 2027 1783 2031 1787 se
tri 2765 1783 2769 1787 sw
rect 2769 1783 2770 1796
rect 2026 1782 2371 1783
rect 2424 1782 2770 1783
rect 2026 1770 2027 1782
tri 2027 1778 2031 1782 ne
tri 2765 1778 2769 1782 nw
rect 2769 1770 2770 1782
rect 3026 1783 3027 1796
tri 3027 1783 3031 1787 se
tri 3765 1783 3769 1787 sw
rect 3769 1783 3770 1796
rect 3026 1782 3371 1783
rect 3424 1782 3770 1783
rect 3026 1770 3027 1782
tri 3027 1778 3031 1782 ne
tri 3765 1778 3769 1782 nw
rect 3769 1770 3770 1782
rect -3847 1620 -3846 1633
tri -3846 1620 -3842 1624 se
tri -3362 1620 -3358 1624 sw
rect -3358 1620 -3357 1633
rect -3847 1619 -3655 1620
rect -3548 1619 -3357 1620
rect -3847 1607 -3846 1619
tri -3846 1615 -3842 1619 ne
tri -3362 1615 -3358 1619 nw
rect -3358 1607 -3357 1619
rect -2847 1620 -2846 1633
tri -2846 1620 -2842 1624 se
tri -2362 1620 -2358 1624 sw
rect -2358 1620 -2357 1633
rect -2847 1619 -2655 1620
rect -2548 1619 -2357 1620
rect -2847 1607 -2846 1619
tri -2846 1615 -2842 1619 ne
tri -2362 1615 -2358 1619 nw
rect -2358 1607 -2357 1619
rect -1847 1620 -1846 1633
tri -1846 1620 -1842 1624 se
tri -1362 1620 -1358 1624 sw
rect -1358 1620 -1357 1633
rect -1847 1619 -1655 1620
rect -1548 1619 -1357 1620
rect -1847 1607 -1846 1619
tri -1846 1615 -1842 1619 ne
tri -1362 1615 -1358 1619 nw
rect -1358 1607 -1357 1619
rect -847 1620 -846 1633
tri -846 1620 -842 1624 se
tri -362 1620 -358 1624 sw
rect -358 1620 -357 1633
rect -847 1619 -655 1620
rect -548 1619 -357 1620
rect -847 1607 -846 1619
tri -846 1615 -842 1619 ne
tri -362 1615 -358 1619 nw
rect -358 1607 -357 1619
rect 153 1620 154 1633
tri 154 1620 158 1624 se
tri 638 1620 642 1624 sw
rect 642 1620 643 1633
rect 153 1619 345 1620
rect 452 1619 643 1620
rect 153 1607 154 1619
tri 154 1615 158 1619 ne
tri 638 1615 642 1619 nw
rect 642 1607 643 1619
rect 1153 1620 1154 1633
tri 1154 1620 1158 1624 se
tri 1638 1620 1642 1624 sw
rect 1642 1620 1643 1633
rect 1153 1619 1345 1620
rect 1452 1619 1643 1620
rect 1153 1607 1154 1619
tri 1154 1615 1158 1619 ne
tri 1638 1615 1642 1619 nw
rect 1642 1607 1643 1619
rect 2153 1620 2154 1633
tri 2154 1620 2158 1624 se
tri 2638 1620 2642 1624 sw
rect 2642 1620 2643 1633
rect 2153 1619 2345 1620
rect 2452 1619 2643 1620
rect 2153 1607 2154 1619
tri 2154 1615 2158 1619 ne
tri 2638 1615 2642 1619 nw
rect 2642 1607 2643 1619
rect 3153 1620 3154 1633
tri 3154 1620 3158 1624 se
tri 3638 1620 3642 1624 sw
rect 3642 1620 3643 1633
rect 3153 1619 3345 1620
rect 3452 1619 3643 1620
rect 3153 1607 3154 1619
tri 3154 1615 3158 1619 ne
tri 3638 1615 3642 1619 nw
rect 3642 1607 3643 1619
rect -3811 1565 -3810 1578
tri -3810 1565 -3806 1569 se
tri -3792 1565 -3788 1569 sw
rect -3788 1565 -3787 1578
rect -3811 1564 -3787 1565
rect -3811 1552 -3810 1564
tri -3810 1560 -3806 1564 ne
tri -3801 1560 -3799 1563 se
tri -3792 1560 -3788 1564 nw
tri -3802 1557 -3801 1560 se
rect -3801 1557 -3799 1560
tri -3799 1557 -3798 1560 sw
rect -3803 1556 -3802 1557
tri -3802 1556 -3801 1557 nw
rect -3799 1556 -3798 1557
rect -3805 1524 -3800 1556
rect -3788 1552 -3787 1564
rect -2811 1565 -2810 1578
tri -2810 1565 -2806 1569 se
tri -2792 1565 -2788 1569 sw
rect -2788 1565 -2787 1578
rect -2811 1564 -2787 1565
rect -2811 1552 -2810 1564
tri -2810 1560 -2806 1564 ne
tri -2801 1560 -2799 1563 se
tri -2792 1560 -2788 1564 nw
tri -2802 1557 -2801 1560 se
rect -2801 1557 -2799 1560
tri -2799 1557 -2798 1560 sw
rect -2803 1556 -2802 1557
tri -2802 1556 -2801 1557 nw
rect -2799 1556 -2798 1557
rect -3393 1533 -3392 1546
tri -3392 1533 -3388 1537 se
tri -3336 1533 -3332 1537 sw
rect -3332 1533 -3331 1546
rect -3393 1532 -3331 1533
rect -3393 1520 -3392 1532
tri -3392 1528 -3388 1532 ne
tri -3336 1528 -3332 1532 nw
rect -3332 1520 -3331 1532
rect -2805 1524 -2800 1556
rect -2788 1552 -2787 1564
rect -1811 1565 -1810 1578
tri -1810 1565 -1806 1569 se
tri -1792 1565 -1788 1569 sw
rect -1788 1565 -1787 1578
rect -1811 1564 -1787 1565
rect -1811 1552 -1810 1564
tri -1810 1560 -1806 1564 ne
tri -1801 1560 -1799 1563 se
tri -1792 1560 -1788 1564 nw
tri -1802 1557 -1801 1560 se
rect -1801 1557 -1799 1560
tri -1799 1557 -1798 1560 sw
rect -1803 1556 -1802 1557
tri -1802 1556 -1801 1557 nw
rect -1799 1556 -1798 1557
rect -2393 1533 -2392 1546
tri -2392 1533 -2388 1537 se
tri -2336 1533 -2332 1537 sw
rect -2332 1533 -2331 1546
rect -2393 1532 -2331 1533
rect -2393 1520 -2392 1532
tri -2392 1528 -2388 1532 ne
tri -2336 1528 -2332 1532 nw
rect -2332 1520 -2331 1532
rect -1805 1524 -1800 1556
rect -1788 1552 -1787 1564
rect -811 1565 -810 1578
tri -810 1565 -806 1569 se
tri -792 1565 -788 1569 sw
rect -788 1565 -787 1578
rect -811 1564 -787 1565
rect -811 1552 -810 1564
tri -810 1560 -806 1564 ne
tri -801 1560 -799 1563 se
tri -792 1560 -788 1564 nw
tri -802 1557 -801 1560 se
rect -801 1557 -799 1560
tri -799 1557 -798 1560 sw
rect -803 1556 -802 1557
tri -802 1556 -801 1557 nw
rect -799 1556 -798 1557
rect -1393 1533 -1392 1546
tri -1392 1533 -1388 1537 se
tri -1336 1533 -1332 1537 sw
rect -1332 1533 -1331 1546
rect -1393 1532 -1331 1533
rect -1393 1520 -1392 1532
tri -1392 1528 -1388 1532 ne
tri -1336 1528 -1332 1532 nw
rect -1332 1520 -1331 1532
rect -805 1524 -800 1556
rect -788 1552 -787 1564
rect 189 1565 190 1578
tri 190 1565 194 1569 se
tri 208 1565 212 1569 sw
rect 212 1565 213 1578
rect 189 1564 213 1565
rect 189 1552 190 1564
tri 190 1560 194 1564 ne
tri 199 1560 201 1563 se
tri 208 1560 212 1564 nw
tri 198 1557 199 1560 se
rect 199 1557 201 1560
tri 201 1557 202 1560 sw
rect 197 1556 198 1557
tri 198 1556 199 1557 nw
rect 201 1556 202 1557
rect -393 1533 -392 1546
tri -392 1533 -388 1537 se
tri -336 1533 -332 1537 sw
rect -332 1533 -331 1546
rect -393 1532 -331 1533
rect -393 1520 -392 1532
tri -392 1528 -388 1532 ne
tri -336 1528 -332 1532 nw
rect -332 1520 -331 1532
rect 195 1524 200 1556
rect 212 1552 213 1564
rect 1189 1565 1190 1578
tri 1190 1565 1194 1569 se
tri 1208 1565 1212 1569 sw
rect 1212 1565 1213 1578
rect 1189 1564 1213 1565
rect 1189 1552 1190 1564
tri 1190 1560 1194 1564 ne
tri 1199 1560 1201 1563 se
tri 1208 1560 1212 1564 nw
tri 1198 1557 1199 1560 se
rect 1199 1557 1201 1560
tri 1201 1557 1202 1560 sw
rect 1197 1556 1198 1557
tri 1198 1556 1199 1557 nw
rect 1201 1556 1202 1557
rect 607 1533 608 1546
tri 608 1533 612 1537 se
tri 664 1533 668 1537 sw
rect 668 1533 669 1546
rect 607 1532 669 1533
rect 607 1520 608 1532
tri 608 1528 612 1532 ne
tri 664 1528 668 1532 nw
rect 668 1520 669 1532
rect 1195 1524 1200 1556
rect 1212 1552 1213 1564
rect 2189 1565 2190 1578
tri 2190 1565 2194 1569 se
tri 2208 1565 2212 1569 sw
rect 2212 1565 2213 1578
rect 2189 1564 2213 1565
rect 2189 1552 2190 1564
tri 2190 1560 2194 1564 ne
tri 2199 1560 2201 1563 se
tri 2208 1560 2212 1564 nw
tri 2198 1557 2199 1560 se
rect 2199 1557 2201 1560
tri 2201 1557 2202 1560 sw
rect 2197 1556 2198 1557
tri 2198 1556 2199 1557 nw
rect 2201 1556 2202 1557
rect 1607 1533 1608 1546
tri 1608 1533 1612 1537 se
tri 1664 1533 1668 1537 sw
rect 1668 1533 1669 1546
rect 1607 1532 1669 1533
rect 1607 1520 1608 1532
tri 1608 1528 1612 1532 ne
tri 1664 1528 1668 1532 nw
rect 1668 1520 1669 1532
rect 2195 1524 2200 1556
rect 2212 1552 2213 1564
rect 3189 1565 3190 1578
tri 3190 1565 3194 1569 se
tri 3208 1565 3212 1569 sw
rect 3212 1565 3213 1578
rect 3189 1564 3213 1565
rect 3189 1552 3190 1564
tri 3190 1560 3194 1564 ne
tri 3199 1560 3201 1563 se
tri 3208 1560 3212 1564 nw
tri 3198 1557 3199 1560 se
rect 3199 1557 3201 1560
tri 3201 1557 3202 1560 sw
rect 3197 1556 3198 1557
tri 3198 1556 3199 1557 nw
rect 3201 1556 3202 1557
rect 2607 1533 2608 1546
tri 2608 1533 2612 1537 se
tri 2664 1533 2668 1537 sw
rect 2668 1533 2669 1546
rect 2607 1532 2669 1533
rect 2607 1520 2608 1532
tri 2608 1528 2612 1532 ne
tri 2664 1528 2668 1532 nw
rect 2668 1520 2669 1532
rect 3195 1524 3200 1556
rect 3212 1552 3213 1564
rect 3607 1533 3608 1546
tri 3608 1533 3612 1537 se
tri 3664 1533 3668 1537 sw
rect 3668 1533 3669 1546
rect 3607 1532 3669 1533
rect 3607 1520 3608 1532
tri 3608 1528 3612 1532 ne
tri 3664 1528 3668 1532 nw
rect 3668 1520 3669 1532
rect -3670 1479 -3669 1492
tri -3669 1479 -3665 1483 se
tri -3539 1479 -3535 1483 sw
rect -3535 1479 -3534 1492
rect -3670 1478 -3623 1479
rect -3581 1478 -3534 1479
rect -3670 1466 -3669 1478
tri -3669 1474 -3665 1478 ne
tri -3539 1474 -3535 1478 nw
rect -3535 1466 -3534 1478
rect -2670 1479 -2669 1492
tri -2669 1479 -2665 1483 se
tri -2539 1479 -2535 1483 sw
rect -2535 1479 -2534 1492
rect -2670 1478 -2623 1479
rect -2581 1478 -2534 1479
rect -2670 1466 -2669 1478
tri -2669 1474 -2665 1478 ne
tri -2539 1474 -2535 1478 nw
rect -2535 1466 -2534 1478
rect -1670 1479 -1669 1492
tri -1669 1479 -1665 1483 se
tri -1539 1479 -1535 1483 sw
rect -1535 1479 -1534 1492
rect -1670 1478 -1623 1479
rect -1581 1478 -1534 1479
rect -1670 1466 -1669 1478
tri -1669 1474 -1665 1478 ne
tri -1539 1474 -1535 1478 nw
rect -1535 1466 -1534 1478
rect -670 1479 -669 1492
tri -669 1479 -665 1483 se
tri -539 1479 -535 1483 sw
rect -535 1479 -534 1492
rect -670 1478 -623 1479
rect -581 1478 -534 1479
rect -670 1466 -669 1478
tri -669 1474 -665 1478 ne
tri -539 1474 -535 1478 nw
rect -535 1466 -534 1478
rect 330 1479 331 1492
tri 331 1479 335 1483 se
tri 461 1479 465 1483 sw
rect 465 1479 466 1492
rect 330 1478 377 1479
rect 419 1478 466 1479
rect 330 1466 331 1478
tri 331 1474 335 1478 ne
tri 461 1474 465 1478 nw
rect 465 1466 466 1478
rect 1330 1479 1331 1492
tri 1331 1479 1335 1483 se
tri 1461 1479 1465 1483 sw
rect 1465 1479 1466 1492
rect 1330 1478 1377 1479
rect 1419 1478 1466 1479
rect 1330 1466 1331 1478
tri 1331 1474 1335 1478 ne
tri 1461 1474 1465 1478 nw
rect 1465 1466 1466 1478
rect 2330 1479 2331 1492
tri 2331 1479 2335 1483 se
tri 2461 1479 2465 1483 sw
rect 2465 1479 2466 1492
rect 2330 1478 2377 1479
rect 2419 1478 2466 1479
rect 2330 1466 2331 1478
tri 2331 1474 2335 1478 ne
tri 2461 1474 2465 1478 nw
rect 2465 1466 2466 1478
rect 3330 1479 3331 1492
tri 3331 1479 3335 1483 se
tri 3461 1479 3465 1483 sw
rect 3465 1479 3466 1492
rect 3330 1478 3377 1479
rect 3419 1478 3466 1479
rect 3330 1466 3331 1478
tri 3331 1474 3335 1478 ne
tri 3461 1474 3465 1478 nw
rect 3465 1466 3466 1478
rect -3811 1442 -3810 1455
tri -3810 1442 -3806 1446 se
tri -3744 1442 -3740 1446 sw
rect -3740 1442 -3739 1455
rect -3811 1441 -3739 1442
rect -3811 1429 -3810 1441
tri -3810 1437 -3806 1441 ne
tri -3744 1437 -3740 1441 nw
rect -3740 1429 -3739 1441
rect -2811 1442 -2810 1455
tri -2810 1442 -2806 1446 se
tri -2744 1442 -2740 1446 sw
rect -2740 1442 -2739 1455
rect -2811 1441 -2739 1442
rect -2811 1429 -2810 1441
tri -2810 1437 -2806 1441 ne
tri -2744 1437 -2740 1441 nw
rect -2740 1429 -2739 1441
rect -1811 1442 -1810 1455
tri -1810 1442 -1806 1446 se
tri -1744 1442 -1740 1446 sw
rect -1740 1442 -1739 1455
rect -1811 1441 -1739 1442
rect -1811 1429 -1810 1441
tri -1810 1437 -1806 1441 ne
tri -1744 1437 -1740 1441 nw
rect -1740 1429 -1739 1441
rect -811 1442 -810 1455
tri -810 1442 -806 1446 se
tri -744 1442 -740 1446 sw
rect -740 1442 -739 1455
rect -811 1441 -739 1442
rect -811 1429 -810 1441
tri -810 1437 -806 1441 ne
tri -744 1437 -740 1441 nw
rect -740 1429 -739 1441
rect 189 1442 190 1455
tri 190 1442 194 1446 se
tri 256 1442 260 1446 sw
rect 260 1442 261 1455
rect 189 1441 261 1442
rect 189 1429 190 1441
tri 190 1437 194 1441 ne
tri 256 1437 260 1441 nw
rect 260 1429 261 1441
rect 1189 1442 1190 1455
tri 1190 1442 1194 1446 se
tri 1256 1442 1260 1446 sw
rect 1260 1442 1261 1455
rect 1189 1441 1261 1442
rect 1189 1429 1190 1441
tri 1190 1437 1194 1441 ne
tri 1256 1437 1260 1441 nw
rect 1260 1429 1261 1441
rect 2189 1442 2190 1455
tri 2190 1442 2194 1446 se
tri 2256 1442 2260 1446 sw
rect 2260 1442 2261 1455
rect 2189 1441 2261 1442
rect 2189 1429 2190 1441
tri 2190 1437 2194 1441 ne
tri 2256 1437 2260 1441 nw
rect 2260 1429 2261 1441
rect 3189 1442 3190 1455
tri 3190 1442 3194 1446 se
tri 3256 1442 3260 1446 sw
rect 3260 1442 3261 1455
rect 3189 1441 3261 1442
rect 3189 1429 3190 1441
tri 3190 1437 3194 1441 ne
tri 3256 1437 3260 1441 nw
rect 3260 1429 3261 1441
tri -3610 1404 -3608 1406 se
tri -3608 1404 -3607 1406 sw
tri -3597 1404 -3596 1406 se
tri -3596 1404 -3594 1406 sw
tri -3610 1403 -3608 1404 ne
rect -3608 1403 -3607 1404
tri -3607 1403 -3605 1404 sw
tri -3599 1403 -3597 1404 se
tri -3608 1400 -3605 1403 ne
tri -3605 1401 -3604 1403 sw
tri -3600 1401 -3599 1403 se
rect -3599 1401 -3597 1403
tri -3597 1401 -3594 1404 nw
tri -2610 1404 -2608 1406 se
tri -2608 1404 -2607 1406 sw
tri -2597 1404 -2596 1406 se
tri -2596 1404 -2594 1406 sw
tri -2610 1403 -2608 1404 ne
rect -2608 1403 -2607 1404
tri -2607 1403 -2605 1404 sw
tri -2599 1403 -2597 1404 se
rect -3605 1400 -3604 1401
tri -3604 1400 -3602 1401 sw
tri -3602 1400 -3600 1401 se
tri -3605 1398 -3604 1400 ne
tri -3607 1395 -3604 1398 se
rect -3604 1396 -3600 1400
tri -3600 1398 -3597 1401 nw
tri -2608 1400 -2605 1403 ne
tri -2605 1401 -2604 1403 sw
tri -2600 1401 -2599 1403 se
rect -2599 1401 -2597 1403
tri -2597 1401 -2594 1404 nw
tri -1610 1404 -1608 1406 se
tri -1608 1404 -1607 1406 sw
tri -1597 1404 -1596 1406 se
tri -1596 1404 -1594 1406 sw
tri -1610 1403 -1608 1404 ne
rect -1608 1403 -1607 1404
tri -1607 1403 -1605 1404 sw
tri -1599 1403 -1597 1404 se
rect -2605 1400 -2604 1401
tri -2604 1400 -2602 1401 sw
tri -2602 1400 -2600 1401 se
tri -2605 1398 -2604 1400 ne
rect -3604 1395 -3603 1396
tri -3603 1395 -3602 1396 nw
tri -3602 1395 -3601 1396 ne
rect -3601 1395 -3600 1396
tri -3600 1395 -3597 1398 sw
tri -2607 1395 -2604 1398 se
rect -2604 1396 -2600 1400
tri -2600 1398 -2597 1401 nw
tri -1608 1400 -1605 1403 ne
tri -1605 1401 -1604 1403 sw
tri -1600 1401 -1599 1403 se
rect -1599 1401 -1597 1403
tri -1597 1401 -1594 1404 nw
tri -610 1404 -608 1406 se
tri -608 1404 -607 1406 sw
tri -597 1404 -596 1406 se
tri -596 1404 -594 1406 sw
tri -610 1403 -608 1404 ne
rect -608 1403 -607 1404
tri -607 1403 -605 1404 sw
tri -599 1403 -597 1404 se
rect -1605 1400 -1604 1401
tri -1604 1400 -1602 1401 sw
tri -1602 1400 -1600 1401 se
tri -1605 1398 -1604 1400 ne
rect -2604 1395 -2603 1396
tri -2603 1395 -2602 1396 nw
tri -2602 1395 -2601 1396 ne
rect -2601 1395 -2600 1396
tri -2600 1395 -2597 1398 sw
tri -1607 1395 -1604 1398 se
rect -1604 1396 -1600 1400
tri -1600 1398 -1597 1401 nw
tri -608 1400 -605 1403 ne
tri -605 1401 -604 1403 sw
tri -600 1401 -599 1403 se
rect -599 1401 -597 1403
tri -597 1401 -594 1404 nw
tri 390 1404 392 1406 se
tri 392 1404 393 1406 sw
tri 403 1404 404 1406 se
tri 404 1404 406 1406 sw
tri 390 1403 392 1404 ne
rect 392 1403 393 1404
tri 393 1403 395 1404 sw
tri 401 1403 403 1404 se
rect -605 1400 -604 1401
tri -604 1400 -602 1401 sw
tri -602 1400 -600 1401 se
tri -605 1398 -604 1400 ne
rect -1604 1395 -1603 1396
tri -1603 1395 -1602 1396 nw
tri -1602 1395 -1601 1396 ne
rect -1601 1395 -1600 1396
tri -1600 1395 -1597 1398 sw
tri -607 1395 -604 1398 se
rect -604 1396 -600 1400
tri -600 1398 -597 1401 nw
tri 392 1400 395 1403 ne
tri 395 1401 396 1403 sw
tri 400 1401 401 1403 se
rect 401 1401 403 1403
tri 403 1401 406 1404 nw
tri 1390 1404 1392 1406 se
tri 1392 1404 1393 1406 sw
tri 1403 1404 1404 1406 se
tri 1404 1404 1406 1406 sw
tri 1390 1403 1392 1404 ne
rect 1392 1403 1393 1404
tri 1393 1403 1395 1404 sw
tri 1401 1403 1403 1404 se
rect 395 1400 396 1401
tri 396 1400 398 1401 sw
tri 398 1400 400 1401 se
tri 395 1398 396 1400 ne
rect -604 1395 -603 1396
tri -603 1395 -602 1396 nw
tri -602 1395 -601 1396 ne
rect -601 1395 -600 1396
tri -600 1395 -597 1398 sw
tri 393 1395 396 1398 se
rect 396 1396 400 1400
tri 400 1398 403 1401 nw
tri 1392 1400 1395 1403 ne
tri 1395 1401 1396 1403 sw
tri 1400 1401 1401 1403 se
rect 1401 1401 1403 1403
tri 1403 1401 1406 1404 nw
tri 2390 1404 2392 1406 se
tri 2392 1404 2393 1406 sw
tri 2403 1404 2404 1406 se
tri 2404 1404 2406 1406 sw
tri 2390 1403 2392 1404 ne
rect 2392 1403 2393 1404
tri 2393 1403 2395 1404 sw
tri 2401 1403 2403 1404 se
rect 1395 1400 1396 1401
tri 1396 1400 1398 1401 sw
tri 1398 1400 1400 1401 se
tri 1395 1398 1396 1400 ne
rect 396 1395 397 1396
tri 397 1395 398 1396 nw
tri 398 1395 399 1396 ne
rect 399 1395 400 1396
tri 400 1395 403 1398 sw
tri 1393 1395 1396 1398 se
rect 1396 1396 1400 1400
tri 1400 1398 1403 1401 nw
tri 2392 1400 2395 1403 ne
tri 2395 1401 2396 1403 sw
tri 2400 1401 2401 1403 se
rect 2401 1401 2403 1403
tri 2403 1401 2406 1404 nw
tri 3390 1404 3392 1406 se
tri 3392 1404 3393 1406 sw
tri 3403 1404 3404 1406 se
tri 3404 1404 3406 1406 sw
tri 3390 1403 3392 1404 ne
rect 3392 1403 3393 1404
tri 3393 1403 3395 1404 sw
tri 3401 1403 3403 1404 se
rect 2395 1400 2396 1401
tri 2396 1400 2398 1401 sw
tri 2398 1400 2400 1401 se
tri 2395 1398 2396 1400 ne
rect 1396 1395 1397 1396
tri 1397 1395 1398 1396 nw
tri 1398 1395 1399 1396 ne
rect 1399 1395 1400 1396
tri 1400 1395 1403 1398 sw
tri 2393 1395 2396 1398 se
rect 2396 1396 2400 1400
tri 2400 1398 2403 1401 nw
tri 3392 1400 3395 1403 ne
tri 3395 1401 3396 1403 sw
tri 3400 1401 3401 1403 se
rect 3401 1401 3403 1403
tri 3403 1401 3406 1404 nw
rect 3395 1400 3396 1401
tri 3396 1400 3398 1401 sw
tri 3398 1400 3400 1401 se
tri 3395 1398 3396 1400 ne
rect 2396 1395 2397 1396
tri 2397 1395 2398 1396 nw
tri 2398 1395 2399 1396 ne
rect 2399 1395 2400 1396
tri 2400 1395 2403 1398 sw
tri 3393 1395 3396 1398 se
rect 3396 1396 3400 1400
tri 3400 1398 3403 1401 nw
rect 3396 1395 3397 1396
tri 3397 1395 3398 1396 nw
tri 3398 1395 3399 1396 ne
rect 3399 1395 3400 1396
tri 3400 1395 3403 1398 sw
tri -3610 1392 -3607 1395 se
tri -3607 1392 -3604 1395 nw
tri -3600 1392 -3597 1395 ne
tri -3597 1392 -3594 1395 sw
tri -3610 1390 -3608 1392 ne
tri -3608 1390 -3607 1392 nw
tri -3597 1390 -3596 1392 ne
tri -3596 1390 -3594 1392 nw
tri -2610 1392 -2607 1395 se
tri -2607 1392 -2604 1395 nw
tri -2600 1392 -2597 1395 ne
tri -2597 1392 -2594 1395 sw
tri -2610 1390 -2608 1392 ne
tri -2608 1390 -2607 1392 nw
tri -2597 1390 -2596 1392 ne
tri -2596 1390 -2594 1392 nw
tri -1610 1392 -1607 1395 se
tri -1607 1392 -1604 1395 nw
tri -1600 1392 -1597 1395 ne
tri -1597 1392 -1594 1395 sw
tri -1610 1390 -1608 1392 ne
tri -1608 1390 -1607 1392 nw
tri -1597 1390 -1596 1392 ne
tri -1596 1390 -1594 1392 nw
tri -610 1392 -607 1395 se
tri -607 1392 -604 1395 nw
tri -600 1392 -597 1395 ne
tri -597 1392 -594 1395 sw
tri -610 1390 -608 1392 ne
tri -608 1390 -607 1392 nw
tri -597 1390 -596 1392 ne
tri -596 1390 -594 1392 nw
tri 390 1392 393 1395 se
tri 393 1392 396 1395 nw
tri 400 1392 403 1395 ne
tri 403 1392 406 1395 sw
tri 390 1390 392 1392 ne
tri 392 1390 393 1392 nw
tri 403 1390 404 1392 ne
tri 404 1390 406 1392 nw
tri 1390 1392 1393 1395 se
tri 1393 1392 1396 1395 nw
tri 1400 1392 1403 1395 ne
tri 1403 1392 1406 1395 sw
tri 1390 1390 1392 1392 ne
tri 1392 1390 1393 1392 nw
tri 1403 1390 1404 1392 ne
tri 1404 1390 1406 1392 nw
tri 2390 1392 2393 1395 se
tri 2393 1392 2396 1395 nw
tri 2400 1392 2403 1395 ne
tri 2403 1392 2406 1395 sw
tri 2390 1390 2392 1392 ne
tri 2392 1390 2393 1392 nw
tri 2403 1390 2404 1392 ne
tri 2404 1390 2406 1392 nw
tri 3390 1392 3393 1395 se
tri 3393 1392 3396 1395 nw
tri 3400 1392 3403 1395 ne
tri 3403 1392 3406 1395 sw
tri 3390 1390 3392 1392 ne
tri 3392 1390 3393 1392 nw
tri 3403 1390 3404 1392 ne
tri 3404 1390 3406 1392 nw
rect -3534 1330 -3533 1343
tri -3533 1330 -3529 1334 se
tri -3470 1330 -3466 1334 sw
rect -3466 1330 -3465 1343
rect -3534 1329 -3465 1330
rect -3534 1317 -3533 1329
tri -3533 1325 -3529 1329 ne
tri -3470 1325 -3466 1329 nw
rect -3466 1317 -3465 1329
rect -3331 1330 -3330 1343
tri -3330 1330 -3326 1334 se
tri -3235 1330 -3231 1334 sw
rect -3231 1330 -3230 1343
rect -3331 1329 -3230 1330
rect -3331 1317 -3330 1329
tri -3330 1325 -3326 1329 ne
tri -3235 1325 -3231 1329 nw
rect -3231 1317 -3230 1329
rect -2534 1330 -2533 1343
tri -2533 1330 -2529 1334 se
tri -2470 1330 -2466 1334 sw
rect -2466 1330 -2465 1343
rect -2534 1329 -2465 1330
rect -2534 1317 -2533 1329
tri -2533 1325 -2529 1329 ne
tri -2470 1325 -2466 1329 nw
rect -2466 1317 -2465 1329
rect -2331 1330 -2330 1343
tri -2330 1330 -2326 1334 se
tri -2235 1330 -2231 1334 sw
rect -2231 1330 -2230 1343
rect -2331 1329 -2230 1330
rect -2331 1317 -2330 1329
tri -2330 1325 -2326 1329 ne
tri -2235 1325 -2231 1329 nw
rect -2231 1317 -2230 1329
rect -1534 1330 -1533 1343
tri -1533 1330 -1529 1334 se
tri -1470 1330 -1466 1334 sw
rect -1466 1330 -1465 1343
rect -1534 1329 -1465 1330
rect -1534 1317 -1533 1329
tri -1533 1325 -1529 1329 ne
tri -1470 1325 -1466 1329 nw
rect -1466 1317 -1465 1329
rect -1331 1330 -1330 1343
tri -1330 1330 -1326 1334 se
tri -1235 1330 -1231 1334 sw
rect -1231 1330 -1230 1343
rect -1331 1329 -1230 1330
rect -1331 1317 -1330 1329
tri -1330 1325 -1326 1329 ne
tri -1235 1325 -1231 1329 nw
rect -1231 1317 -1230 1329
rect -534 1330 -533 1343
tri -533 1330 -529 1334 se
tri -470 1330 -466 1334 sw
rect -466 1330 -465 1343
rect -534 1329 -465 1330
rect -534 1317 -533 1329
tri -533 1325 -529 1329 ne
tri -470 1325 -466 1329 nw
rect -466 1317 -465 1329
rect -331 1330 -330 1343
tri -330 1330 -326 1334 se
tri -235 1330 -231 1334 sw
rect -231 1330 -230 1343
rect -331 1329 -230 1330
rect -331 1317 -330 1329
tri -330 1325 -326 1329 ne
tri -235 1325 -231 1329 nw
rect -231 1317 -230 1329
rect 466 1330 467 1343
tri 467 1330 471 1334 se
tri 530 1330 534 1334 sw
rect 534 1330 535 1343
rect 466 1329 535 1330
rect 466 1317 467 1329
tri 467 1325 471 1329 ne
tri 530 1325 534 1329 nw
rect 534 1317 535 1329
rect 669 1330 670 1343
tri 670 1330 674 1334 se
tri 765 1330 769 1334 sw
rect 769 1330 770 1343
rect 669 1329 770 1330
rect 669 1317 670 1329
tri 670 1325 674 1329 ne
tri 765 1325 769 1329 nw
rect 769 1317 770 1329
rect 1466 1330 1467 1343
tri 1467 1330 1471 1334 se
tri 1530 1330 1534 1334 sw
rect 1534 1330 1535 1343
rect 1466 1329 1535 1330
rect 1466 1317 1467 1329
tri 1467 1325 1471 1329 ne
tri 1530 1325 1534 1329 nw
rect 1534 1317 1535 1329
rect 1669 1330 1670 1343
tri 1670 1330 1674 1334 se
tri 1765 1330 1769 1334 sw
rect 1769 1330 1770 1343
rect 1669 1329 1770 1330
rect 1669 1317 1670 1329
tri 1670 1325 1674 1329 ne
tri 1765 1325 1769 1329 nw
rect 1769 1317 1770 1329
rect 2466 1330 2467 1343
tri 2467 1330 2471 1334 se
tri 2530 1330 2534 1334 sw
rect 2534 1330 2535 1343
rect 2466 1329 2535 1330
rect 2466 1317 2467 1329
tri 2467 1325 2471 1329 ne
tri 2530 1325 2534 1329 nw
rect 2534 1317 2535 1329
rect 2669 1330 2670 1343
tri 2670 1330 2674 1334 se
tri 2765 1330 2769 1334 sw
rect 2769 1330 2770 1343
rect 2669 1329 2770 1330
rect 2669 1317 2670 1329
tri 2670 1325 2674 1329 ne
tri 2765 1325 2769 1329 nw
rect 2769 1317 2770 1329
rect 3466 1330 3467 1343
tri 3467 1330 3471 1334 se
tri 3530 1330 3534 1334 sw
rect 3534 1330 3535 1343
rect 3466 1329 3535 1330
rect 3466 1317 3467 1329
tri 3467 1325 3471 1329 ne
tri 3530 1325 3534 1329 nw
rect 3534 1317 3535 1329
rect 3669 1330 3670 1343
tri 3670 1330 3674 1334 se
tri 3765 1330 3769 1334 sw
rect 3769 1330 3770 1343
rect 3669 1329 3770 1330
rect 3669 1317 3670 1329
tri 3670 1325 3674 1329 ne
tri 3765 1325 3769 1329 nw
rect 3769 1317 3770 1329
rect -3811 1176 -3810 1189
tri -3810 1176 -3806 1180 se
tri -3398 1176 -3394 1180 sw
rect -3394 1176 -3393 1189
rect -3811 1175 -3623 1176
rect -3581 1175 -3393 1176
rect -3811 1163 -3810 1175
tri -3810 1171 -3806 1175 ne
tri -3398 1171 -3394 1175 nw
rect -3394 1163 -3393 1175
rect -2811 1176 -2810 1189
tri -2810 1176 -2806 1180 se
tri -2398 1176 -2394 1180 sw
rect -2394 1176 -2393 1189
rect -2811 1175 -2623 1176
rect -2581 1175 -2393 1176
rect -2811 1163 -2810 1175
tri -2810 1171 -2806 1175 ne
tri -2398 1171 -2394 1175 nw
rect -2394 1163 -2393 1175
rect -1811 1176 -1810 1189
tri -1810 1176 -1806 1180 se
tri -1398 1176 -1394 1180 sw
rect -1394 1176 -1393 1189
rect -1811 1175 -1623 1176
rect -1581 1175 -1393 1176
rect -1811 1163 -1810 1175
tri -1810 1171 -1806 1175 ne
tri -1398 1171 -1394 1175 nw
rect -1394 1163 -1393 1175
rect -811 1176 -810 1189
tri -810 1176 -806 1180 se
tri -398 1176 -394 1180 sw
rect -394 1176 -393 1189
rect -811 1175 -623 1176
rect -581 1175 -393 1176
rect -811 1163 -810 1175
tri -810 1171 -806 1175 ne
tri -398 1171 -394 1175 nw
rect -394 1163 -393 1175
rect 189 1176 190 1189
tri 190 1176 194 1180 se
tri 602 1176 606 1180 sw
rect 606 1176 607 1189
rect 189 1175 377 1176
rect 419 1175 607 1176
rect 189 1163 190 1175
tri 190 1171 194 1175 ne
tri 602 1171 606 1175 nw
rect 606 1163 607 1175
rect 1189 1176 1190 1189
tri 1190 1176 1194 1180 se
tri 1602 1176 1606 1180 sw
rect 1606 1176 1607 1189
rect 1189 1175 1377 1176
rect 1419 1175 1607 1176
rect 1189 1163 1190 1175
tri 1190 1171 1194 1175 ne
tri 1602 1171 1606 1175 nw
rect 1606 1163 1607 1175
rect 2189 1176 2190 1189
tri 2190 1176 2194 1180 se
tri 2602 1176 2606 1180 sw
rect 2606 1176 2607 1189
rect 2189 1175 2377 1176
rect 2419 1175 2607 1176
rect 2189 1163 2190 1175
tri 2190 1171 2194 1175 ne
tri 2602 1171 2606 1175 nw
rect 2606 1163 2607 1175
rect 3189 1176 3190 1189
tri 3190 1176 3194 1180 se
tri 3602 1176 3606 1180 sw
rect 3606 1176 3607 1189
rect 3189 1175 3377 1176
rect 3419 1175 3607 1176
rect 3189 1163 3190 1175
tri 3190 1171 3194 1175 ne
tri 3602 1171 3606 1175 nw
rect 3606 1163 3607 1175
rect -3638 1136 -3637 1149
tri -3637 1136 -3633 1140 se
tri -3571 1136 -3567 1140 sw
rect -3567 1136 -3566 1149
rect -3638 1135 -3566 1136
rect -3638 1123 -3637 1135
tri -3637 1131 -3633 1135 ne
tri -3571 1131 -3567 1135 nw
rect -3567 1123 -3566 1135
rect -2638 1136 -2637 1149
tri -2637 1136 -2633 1140 se
tri -2571 1136 -2567 1140 sw
rect -2567 1136 -2566 1149
rect -2638 1135 -2566 1136
rect -2638 1123 -2637 1135
tri -2637 1131 -2633 1135 ne
tri -2571 1131 -2567 1135 nw
rect -2567 1123 -2566 1135
rect -1638 1136 -1637 1149
tri -1637 1136 -1633 1140 se
tri -1571 1136 -1567 1140 sw
rect -1567 1136 -1566 1149
rect -1638 1135 -1566 1136
rect -1638 1123 -1637 1135
tri -1637 1131 -1633 1135 ne
tri -1571 1131 -1567 1135 nw
rect -1567 1123 -1566 1135
rect -638 1136 -637 1149
tri -637 1136 -633 1140 se
tri -571 1136 -567 1140 sw
rect -567 1136 -566 1149
rect -638 1135 -566 1136
rect -638 1123 -637 1135
tri -637 1131 -633 1135 ne
tri -571 1131 -567 1135 nw
rect -567 1123 -566 1135
rect 362 1136 363 1149
tri 363 1136 367 1140 se
tri 429 1136 433 1140 sw
rect 433 1136 434 1149
rect 362 1135 434 1136
rect 362 1123 363 1135
tri 363 1131 367 1135 ne
tri 429 1131 433 1135 nw
rect 433 1123 434 1135
rect 1362 1136 1363 1149
tri 1363 1136 1367 1140 se
tri 1429 1136 1433 1140 sw
rect 1433 1136 1434 1149
rect 1362 1135 1434 1136
rect 1362 1123 1363 1135
tri 1363 1131 1367 1135 ne
tri 1429 1131 1433 1135 nw
rect 1433 1123 1434 1135
rect 2362 1136 2363 1149
tri 2363 1136 2367 1140 se
tri 2429 1136 2433 1140 sw
rect 2433 1136 2434 1149
rect 2362 1135 2434 1136
rect 2362 1123 2363 1135
tri 2363 1131 2367 1135 ne
tri 2429 1131 2433 1135 nw
rect 2433 1123 2434 1135
rect 3362 1136 3363 1149
tri 3363 1136 3367 1140 se
tri 3429 1136 3433 1140 sw
rect 3433 1136 3434 1149
rect 3362 1135 3434 1136
rect 3362 1123 3363 1135
tri 3363 1131 3367 1135 ne
tri 3429 1131 3433 1135 nw
rect 3433 1123 3434 1135
rect -3974 783 -3973 796
tri -3973 783 -3969 787 se
tri -3235 783 -3231 787 sw
rect -3231 783 -3230 796
rect -3974 782 -3629 783
rect -3576 782 -3230 783
rect -3974 770 -3973 782
tri -3973 778 -3969 782 ne
tri -3235 778 -3231 782 nw
rect -3231 770 -3230 782
rect -2974 783 -2973 796
tri -2973 783 -2969 787 se
tri -2235 783 -2231 787 sw
rect -2231 783 -2230 796
rect -2974 782 -2629 783
rect -2576 782 -2230 783
rect -2974 770 -2973 782
tri -2973 778 -2969 782 ne
tri -2235 778 -2231 782 nw
rect -2231 770 -2230 782
rect -1974 783 -1973 796
tri -1973 783 -1969 787 se
tri -1235 783 -1231 787 sw
rect -1231 783 -1230 796
rect -1974 782 -1629 783
rect -1576 782 -1230 783
rect -1974 770 -1973 782
tri -1973 778 -1969 782 ne
tri -1235 778 -1231 782 nw
rect -1231 770 -1230 782
rect -974 783 -973 796
tri -973 783 -969 787 se
tri -235 783 -231 787 sw
rect -231 783 -230 796
rect -974 782 -629 783
rect -576 782 -230 783
rect -974 770 -973 782
tri -973 778 -969 782 ne
tri -235 778 -231 782 nw
rect -231 770 -230 782
rect 1026 783 1027 796
tri 1027 783 1031 787 se
tri 1765 783 1769 787 sw
rect 1769 783 1770 796
rect 1026 782 1371 783
rect 1424 782 1770 783
rect 1026 770 1027 782
tri 1027 778 1031 782 ne
tri 1765 778 1769 782 nw
rect 1769 770 1770 782
rect 2026 783 2027 796
tri 2027 783 2031 787 se
tri 2765 783 2769 787 sw
rect 2769 783 2770 796
rect 2026 782 2371 783
rect 2424 782 2770 783
rect 2026 770 2027 782
tri 2027 778 2031 782 ne
tri 2765 778 2769 782 nw
rect 2769 770 2770 782
rect 3026 783 3027 796
tri 3027 783 3031 787 se
tri 3765 783 3769 787 sw
rect 3769 783 3770 796
rect 3026 782 3371 783
rect 3424 782 3770 783
rect 3026 770 3027 782
tri 3027 778 3031 782 ne
tri 3765 778 3769 782 nw
rect 3769 770 3770 782
rect -3847 620 -3846 633
tri -3846 620 -3842 624 se
tri -3362 620 -3358 624 sw
rect -3358 620 -3357 633
rect -3847 619 -3655 620
rect -3548 619 -3357 620
rect -3847 607 -3846 619
tri -3846 615 -3842 619 ne
tri -3362 615 -3358 619 nw
rect -3358 607 -3357 619
rect -2847 620 -2846 633
tri -2846 620 -2842 624 se
tri -2362 620 -2358 624 sw
rect -2358 620 -2357 633
rect -2847 619 -2655 620
rect -2548 619 -2357 620
rect -2847 607 -2846 619
tri -2846 615 -2842 619 ne
tri -2362 615 -2358 619 nw
rect -2358 607 -2357 619
rect -1847 620 -1846 633
tri -1846 620 -1842 624 se
tri -1362 620 -1358 624 sw
rect -1358 620 -1357 633
rect -1847 619 -1655 620
rect -1548 619 -1357 620
rect -1847 607 -1846 619
tri -1846 615 -1842 619 ne
tri -1362 615 -1358 619 nw
rect -1358 607 -1357 619
rect -847 620 -846 633
tri -846 620 -842 624 se
tri -362 620 -358 624 sw
rect -358 620 -357 633
rect -847 619 -655 620
rect -548 619 -357 620
rect -847 607 -846 619
tri -846 615 -842 619 ne
tri -362 615 -358 619 nw
rect -358 607 -357 619
rect 1153 620 1154 633
tri 1154 620 1158 624 se
tri 1638 620 1642 624 sw
rect 1642 620 1643 633
rect 1153 619 1345 620
rect 1452 619 1643 620
rect 1153 607 1154 619
tri 1154 615 1158 619 ne
tri 1638 615 1642 619 nw
rect 1642 607 1643 619
rect 2153 620 2154 633
tri 2154 620 2158 624 se
tri 2638 620 2642 624 sw
rect 2642 620 2643 633
rect 2153 619 2345 620
rect 2452 619 2643 620
rect 2153 607 2154 619
tri 2154 615 2158 619 ne
tri 2638 615 2642 619 nw
rect 2642 607 2643 619
rect 3153 620 3154 633
tri 3154 620 3158 624 se
tri 3638 620 3642 624 sw
rect 3642 620 3643 633
rect 3153 619 3345 620
rect 3452 619 3643 620
rect 3153 607 3154 619
tri 3154 615 3158 619 ne
tri 3638 615 3642 619 nw
rect 3642 607 3643 619
rect -3811 565 -3810 578
tri -3810 565 -3806 569 se
tri -3792 565 -3788 569 sw
rect -3788 565 -3787 578
rect -3811 564 -3787 565
rect -3811 552 -3810 564
tri -3810 560 -3806 564 ne
tri -3801 560 -3799 563 se
tri -3792 560 -3788 564 nw
tri -3802 557 -3801 560 se
rect -3801 557 -3799 560
tri -3799 557 -3798 560 sw
rect -3803 556 -3802 557
tri -3802 556 -3801 557 nw
rect -3799 556 -3798 557
rect -3805 524 -3800 556
rect -3788 552 -3787 564
rect -2811 565 -2810 578
tri -2810 565 -2806 569 se
tri -2792 565 -2788 569 sw
rect -2788 565 -2787 578
rect -2811 564 -2787 565
rect -2811 552 -2810 564
tri -2810 560 -2806 564 ne
tri -2801 560 -2799 563 se
tri -2802 557 -2801 560 se
rect -2801 557 -2799 560
tri -2799 557 -2798 563 sw
tri -2792 560 -2788 564 nw
rect -2803 556 -2802 557
tri -2802 556 -2801 557 nw
rect -2799 556 -2798 557
rect -3393 533 -3392 546
tri -3392 533 -3388 537 se
tri -3336 533 -3332 537 sw
rect -3332 533 -3331 546
rect -3393 532 -3331 533
rect -3393 520 -3392 532
tri -3392 528 -3388 532 ne
tri -3336 528 -3332 532 nw
rect -3332 520 -3331 532
rect -2805 524 -2800 556
rect -2788 552 -2787 564
rect -1811 565 -1810 578
tri -1810 565 -1806 569 se
tri -1792 565 -1788 569 sw
rect -1788 565 -1787 578
rect -1811 564 -1787 565
rect -1811 552 -1810 564
tri -1810 560 -1806 564 ne
tri -1801 560 -1799 563 se
tri -1792 560 -1788 564 nw
tri -1802 557 -1801 560 se
rect -1801 557 -1799 560
tri -1799 557 -1798 560 sw
rect -1803 556 -1802 557
tri -1802 556 -1801 557 nw
rect -1799 556 -1798 557
rect -2393 533 -2392 546
tri -2392 533 -2388 537 se
tri -2336 533 -2332 537 sw
rect -2332 533 -2331 546
rect -2393 532 -2331 533
rect -2393 520 -2392 532
tri -2392 528 -2388 532 ne
tri -2336 528 -2332 532 nw
rect -2332 520 -2331 532
rect -1805 524 -1800 556
rect -1788 552 -1787 564
rect -811 565 -810 578
tri -810 565 -806 569 se
tri -792 565 -788 569 sw
rect -788 565 -787 578
rect -811 564 -787 565
rect -811 552 -810 564
tri -810 560 -806 564 ne
tri -801 560 -799 563 se
tri -792 560 -788 564 nw
tri -802 557 -801 560 se
rect -801 557 -799 560
tri -799 557 -798 560 sw
rect -803 556 -802 557
tri -802 556 -801 557 nw
rect -799 556 -798 557
rect -1393 533 -1392 546
tri -1392 533 -1388 537 se
tri -1336 533 -1332 537 sw
rect -1332 533 -1331 546
rect -1393 532 -1331 533
rect -1393 520 -1392 532
tri -1392 528 -1388 532 ne
tri -1336 528 -1332 532 nw
rect -1332 520 -1331 532
rect -805 524 -800 556
rect -788 552 -787 564
rect 1189 565 1190 578
tri 1190 565 1194 569 se
tri 1208 565 1212 569 sw
rect 1212 565 1213 578
rect 1189 564 1213 565
rect 1189 552 1190 564
tri 1190 560 1194 564 ne
tri 1199 560 1201 563 se
tri 1208 560 1212 564 nw
tri 1198 557 1199 560 se
rect 1199 557 1201 560
tri 1201 557 1202 560 sw
rect 1197 556 1198 557
tri 1198 556 1199 557 nw
rect 1201 556 1202 557
rect -393 533 -392 546
tri -392 533 -388 537 se
tri -336 533 -332 537 sw
rect -332 533 -331 546
rect -393 532 -331 533
rect -393 520 -392 532
tri -392 528 -388 532 ne
tri -336 528 -332 532 nw
rect -332 520 -331 532
rect 1195 524 1200 556
rect 1212 552 1213 564
rect 2189 565 2190 578
tri 2190 565 2194 569 se
tri 2208 565 2212 569 sw
rect 2212 565 2213 578
rect 2189 564 2213 565
rect 2189 552 2190 564
tri 2190 560 2194 564 ne
tri 2199 560 2201 563 se
tri 2208 560 2212 564 nw
tri 2198 557 2199 560 se
rect 2199 557 2201 560
tri 2201 557 2202 560 sw
rect 2197 556 2198 557
tri 2198 556 2199 557 nw
rect 2201 556 2202 557
rect 1607 533 1608 546
tri 1608 533 1612 537 se
tri 1664 533 1668 537 sw
rect 1668 533 1669 546
rect 1607 532 1669 533
rect 1607 520 1608 532
tri 1608 528 1612 532 ne
tri 1664 528 1668 532 nw
rect 1668 520 1669 532
rect 2195 524 2200 556
rect 2212 552 2213 564
rect 3189 565 3190 578
tri 3190 565 3194 569 se
tri 3208 565 3212 569 sw
rect 3212 565 3213 578
rect 3189 564 3213 565
rect 3189 552 3190 564
tri 3190 560 3194 564 ne
tri 3199 560 3201 563 se
tri 3208 560 3212 564 nw
tri 3198 557 3199 560 se
rect 3199 557 3201 560
tri 3201 557 3202 560 sw
rect 3197 556 3198 557
tri 3198 556 3199 557 nw
rect 3201 556 3202 557
rect 2607 533 2608 546
tri 2608 533 2612 537 se
tri 2664 533 2668 537 sw
rect 2668 533 2669 546
rect 2607 532 2669 533
rect 2607 520 2608 532
tri 2608 528 2612 532 ne
tri 2664 528 2668 532 nw
rect 2668 520 2669 532
rect 3195 524 3200 556
rect 3212 552 3213 564
rect 3607 533 3608 546
tri 3608 533 3612 537 se
tri 3664 533 3668 537 sw
rect 3668 533 3669 546
rect 3607 532 3669 533
rect 3607 520 3608 532
tri 3608 528 3612 532 ne
tri 3664 528 3668 532 nw
rect 3668 520 3669 532
rect -3670 479 -3669 492
tri -3669 479 -3665 483 se
tri -3539 479 -3535 483 sw
rect -3535 479 -3534 492
rect -3670 478 -3623 479
rect -3581 478 -3534 479
rect -3670 466 -3669 478
tri -3669 474 -3665 478 ne
tri -3539 474 -3535 478 nw
rect -3535 466 -3534 478
rect -2670 479 -2669 492
tri -2669 479 -2665 483 se
tri -2539 479 -2535 483 sw
rect -2535 479 -2534 492
rect -2670 478 -2623 479
rect -2581 478 -2534 479
rect -2670 466 -2669 478
tri -2669 474 -2665 478 ne
tri -2539 474 -2535 478 nw
rect -2535 466 -2534 478
rect -1670 479 -1669 492
tri -1669 479 -1665 483 se
tri -1539 479 -1535 483 sw
rect -1535 479 -1534 492
rect -1670 478 -1623 479
rect -1581 478 -1534 479
rect -1670 466 -1669 478
tri -1669 474 -1665 478 ne
tri -1539 474 -1535 478 nw
rect -1535 466 -1534 478
rect -670 479 -669 492
tri -669 479 -665 483 se
tri -539 479 -535 483 sw
rect -535 479 -534 492
rect -670 478 -623 479
rect -581 478 -534 479
rect -670 466 -669 478
tri -669 474 -665 478 ne
tri -539 474 -535 478 nw
rect -535 466 -534 478
rect 1330 479 1331 492
tri 1331 479 1335 483 se
tri 1461 479 1465 483 sw
rect 1465 479 1466 492
rect 1330 478 1377 479
rect 1419 478 1466 479
rect 1330 466 1331 478
tri 1331 474 1335 478 ne
tri 1461 474 1465 478 nw
rect 1465 466 1466 478
rect 2330 479 2331 492
tri 2331 479 2335 483 se
tri 2461 479 2465 483 sw
rect 2465 479 2466 492
rect 2330 478 2377 479
rect 2419 478 2466 479
rect 2330 466 2331 478
tri 2331 474 2335 478 ne
tri 2461 474 2465 478 nw
rect 2465 466 2466 478
rect 3330 479 3331 492
tri 3331 479 3335 483 se
tri 3461 479 3465 483 sw
rect 3465 479 3466 492
rect 3330 478 3377 479
rect 3419 478 3466 479
rect 3330 466 3331 478
tri 3331 474 3335 478 ne
tri 3461 474 3465 478 nw
rect 3465 466 3466 478
rect -3811 442 -3810 455
tri -3810 442 -3806 446 se
tri -3744 442 -3740 446 sw
rect -3740 442 -3739 455
rect -3811 441 -3739 442
rect -3811 429 -3810 441
tri -3810 437 -3806 441 ne
tri -3744 437 -3740 441 nw
rect -3740 429 -3739 441
rect -2811 442 -2810 455
tri -2810 442 -2806 446 se
tri -2744 442 -2740 446 sw
rect -2740 442 -2739 455
rect -2811 441 -2739 442
rect -2811 429 -2810 441
tri -2810 437 -2806 441 ne
tri -2744 437 -2740 441 nw
rect -2740 429 -2739 441
rect -1811 442 -1810 455
tri -1810 442 -1806 446 se
tri -1744 442 -1740 446 sw
rect -1740 442 -1739 455
rect -1811 441 -1739 442
rect -1811 429 -1810 441
tri -1810 437 -1806 441 ne
tri -1744 437 -1740 441 nw
rect -1740 429 -1739 441
rect -811 442 -810 455
tri -810 442 -806 446 se
tri -744 442 -740 446 sw
rect -740 442 -739 455
rect -811 441 -739 442
rect -811 429 -810 441
tri -810 437 -806 441 ne
tri -744 437 -740 441 nw
rect -740 429 -739 441
rect 1189 442 1190 455
tri 1190 442 1194 446 se
tri 1256 442 1260 446 sw
rect 1260 442 1261 455
rect 1189 441 1261 442
rect 1189 429 1190 441
tri 1190 437 1194 441 ne
tri 1256 437 1260 441 nw
rect 1260 429 1261 441
rect 2189 442 2190 455
tri 2190 442 2194 446 se
tri 2256 442 2260 446 sw
rect 2260 442 2261 455
rect 2189 441 2261 442
rect 2189 429 2190 441
tri 2190 437 2194 441 ne
tri 2256 437 2260 441 nw
rect 2260 429 2261 441
rect 3189 442 3190 455
tri 3190 442 3194 446 se
tri 3256 442 3260 446 sw
rect 3260 442 3261 455
rect 3189 441 3261 442
rect 3189 429 3190 441
tri 3190 437 3194 441 ne
tri 3256 437 3260 441 nw
rect 3260 429 3261 441
tri -3610 404 -3608 406 se
tri -3608 404 -3607 406 sw
tri -3597 404 -3596 406 se
tri -3596 404 -3594 406 sw
tri -3610 403 -3608 404 ne
rect -3608 403 -3607 404
tri -3607 403 -3605 404 sw
tri -3599 403 -3597 404 se
tri -3608 400 -3605 403 ne
tri -3605 401 -3604 403 sw
tri -3600 401 -3599 403 se
rect -3599 401 -3597 403
tri -3597 401 -3594 404 nw
tri -2610 404 -2608 406 se
tri -2608 404 -2607 406 sw
tri -2597 404 -2596 406 se
tri -2596 404 -2594 406 sw
tri -2610 403 -2608 404 ne
rect -2608 403 -2607 404
tri -2607 403 -2605 404 sw
tri -2599 403 -2597 404 se
rect -3605 400 -3604 401
tri -3604 400 -3602 401 sw
tri -3602 400 -3600 401 se
tri -3605 398 -3604 400 ne
tri -3607 395 -3604 398 se
rect -3604 396 -3600 400
tri -3600 398 -3597 401 nw
tri -2608 400 -2605 403 ne
tri -2605 401 -2604 403 sw
tri -2600 401 -2599 403 se
rect -2599 401 -2597 403
tri -2597 401 -2594 404 nw
tri -1610 404 -1608 406 se
tri -1608 404 -1607 406 sw
tri -1597 404 -1596 406 se
tri -1596 404 -1594 406 sw
tri -1610 403 -1608 404 ne
rect -1608 403 -1607 404
tri -1607 403 -1605 404 sw
tri -1599 403 -1597 404 se
rect -2605 400 -2604 401
tri -2604 400 -2602 401 sw
tri -2602 400 -2600 401 se
tri -2605 398 -2604 400 ne
rect -3604 395 -3603 396
tri -3603 395 -3602 396 nw
tri -3602 395 -3601 396 ne
rect -3601 395 -3600 396
tri -3600 395 -3597 398 sw
tri -2607 395 -2604 398 se
rect -2604 396 -2600 400
tri -2600 398 -2597 401 nw
tri -1608 400 -1605 403 ne
tri -1605 401 -1604 403 sw
tri -1600 401 -1599 403 se
rect -1599 401 -1597 403
tri -1597 401 -1594 404 nw
tri -610 404 -608 406 se
tri -608 404 -607 406 sw
tri -597 404 -596 406 se
tri -596 404 -594 406 sw
tri -610 403 -608 404 ne
rect -608 403 -607 404
tri -607 403 -605 404 sw
tri -599 403 -597 404 se
rect -1605 400 -1604 401
tri -1604 400 -1602 401 sw
tri -1602 400 -1600 401 se
tri -1605 398 -1604 400 ne
rect -2604 395 -2603 396
tri -2603 395 -2602 396 nw
tri -2602 395 -2601 396 ne
rect -2601 395 -2600 396
tri -2600 395 -2597 398 sw
tri -1607 395 -1604 398 se
rect -1604 396 -1600 400
tri -1600 398 -1597 401 nw
tri -608 400 -605 403 ne
tri -605 401 -604 403 sw
tri -600 401 -599 403 se
rect -599 401 -597 403
tri -597 401 -594 404 nw
tri 1390 404 1392 406 se
tri 1392 404 1393 406 sw
tri 1403 404 1404 406 se
tri 1404 404 1406 406 sw
tri 1390 403 1392 404 ne
rect 1392 403 1393 404
tri 1393 403 1395 404 sw
tri 1401 403 1403 404 se
rect -605 400 -604 401
tri -604 400 -602 401 sw
tri -602 400 -600 401 se
tri -605 398 -604 400 ne
rect -1604 395 -1603 396
tri -1603 395 -1602 396 nw
tri -1602 395 -1601 396 ne
rect -1601 395 -1600 396
tri -1600 395 -1597 398 sw
tri -607 395 -604 398 se
rect -604 396 -600 400
tri -600 398 -597 401 nw
tri 1392 400 1395 403 ne
tri 1395 401 1396 403 sw
tri 1400 401 1401 403 se
rect 1401 401 1403 403
tri 1403 401 1406 404 nw
tri 2390 404 2392 406 se
tri 2392 404 2393 406 sw
tri 2403 404 2404 406 se
tri 2404 404 2406 406 sw
tri 2390 403 2392 404 ne
rect 2392 403 2393 404
tri 2393 403 2395 404 sw
tri 2401 403 2403 404 se
rect 1395 400 1396 401
tri 1396 400 1398 401 sw
tri 1398 400 1400 401 se
tri 1395 398 1396 400 ne
rect -604 395 -603 396
tri -603 395 -602 396 nw
tri -602 395 -601 396 ne
rect -601 395 -600 396
tri -600 395 -597 398 sw
tri 1393 395 1396 398 se
rect 1396 396 1400 400
tri 1400 398 1403 401 nw
tri 2392 400 2395 403 ne
tri 2395 401 2396 403 sw
tri 2400 401 2401 403 se
rect 2401 401 2403 403
tri 2403 401 2406 404 nw
tri 3390 404 3392 406 se
tri 3392 404 3393 406 sw
tri 3403 404 3404 406 se
tri 3404 404 3406 406 sw
tri 3390 403 3392 404 ne
rect 3392 403 3393 404
tri 3393 403 3395 404 sw
tri 3401 403 3403 404 se
rect 2395 400 2396 401
tri 2396 400 2398 401 sw
tri 2398 400 2400 401 se
tri 2395 398 2396 400 ne
rect 1396 395 1397 396
tri 1397 395 1398 396 nw
tri 1398 395 1399 396 ne
rect 1399 395 1400 396
tri 1400 395 1403 398 sw
tri 2393 395 2396 398 se
rect 2396 396 2400 400
tri 2400 398 2403 401 nw
tri 3392 400 3395 403 ne
tri 3395 401 3396 403 sw
tri 3400 401 3401 403 se
rect 3401 401 3403 403
tri 3403 401 3406 404 nw
rect 3395 400 3396 401
tri 3396 400 3398 401 sw
tri 3398 400 3400 401 se
tri 3395 398 3396 400 ne
rect 2396 395 2397 396
tri 2397 395 2398 396 nw
tri 2398 395 2399 396 ne
rect 2399 395 2400 396
tri 2400 395 2403 398 sw
tri 3393 395 3396 398 se
rect 3396 396 3400 400
tri 3400 398 3403 401 nw
rect 3396 395 3397 396
tri 3397 395 3398 396 nw
tri 3398 395 3399 396 ne
rect 3399 395 3400 396
tri 3400 395 3403 398 sw
tri -3610 392 -3607 395 se
tri -3607 392 -3604 395 nw
tri -3600 392 -3597 395 ne
tri -3597 392 -3594 395 sw
tri -3610 390 -3608 392 ne
tri -3608 390 -3607 392 nw
tri -3597 390 -3596 392 ne
tri -3596 390 -3594 392 nw
tri -2610 392 -2607 395 se
tri -2607 392 -2604 395 nw
tri -2600 392 -2597 395 ne
tri -2597 392 -2594 395 sw
tri -2610 390 -2608 392 ne
tri -2608 390 -2607 392 nw
tri -2597 390 -2596 392 ne
tri -2596 390 -2594 392 nw
tri -1610 392 -1607 395 se
tri -1607 392 -1604 395 nw
tri -1600 392 -1597 395 ne
tri -1597 392 -1594 395 sw
tri -1610 390 -1608 392 ne
tri -1608 390 -1607 392 nw
tri -1597 390 -1596 392 ne
tri -1596 390 -1594 392 nw
tri -610 392 -607 395 se
tri -607 392 -604 395 nw
tri -600 392 -597 395 ne
tri -597 392 -594 395 sw
tri -610 390 -608 392 ne
tri -608 390 -607 392 nw
tri -597 390 -596 392 ne
tri -596 390 -594 392 nw
tri 1390 392 1393 395 se
tri 1393 392 1396 395 nw
tri 1400 392 1403 395 ne
tri 1403 392 1406 395 sw
tri 1390 390 1392 392 ne
tri 1392 390 1393 392 nw
tri 1403 390 1404 392 ne
tri 1404 390 1406 392 nw
tri 2390 392 2393 395 se
tri 2393 392 2396 395 nw
tri 2400 392 2403 395 ne
tri 2403 392 2406 395 sw
tri 2390 390 2392 392 ne
tri 2392 390 2393 392 nw
tri 2403 390 2404 392 ne
tri 2404 390 2406 392 nw
tri 3390 392 3393 395 se
tri 3393 392 3396 395 nw
tri 3400 392 3403 395 ne
tri 3403 392 3406 395 sw
tri 3390 390 3392 392 ne
tri 3392 390 3393 392 nw
tri 3403 390 3404 392 ne
tri 3404 390 3406 392 nw
rect -3534 330 -3533 343
tri -3533 330 -3529 334 se
tri -3470 330 -3466 334 sw
rect -3466 330 -3465 343
rect -3534 329 -3465 330
rect -3534 317 -3533 329
tri -3533 325 -3529 329 ne
tri -3470 325 -3466 329 nw
rect -3466 317 -3465 329
rect -3331 330 -3330 343
tri -3330 330 -3326 334 se
tri -3235 330 -3231 334 sw
rect -3231 330 -3230 343
rect -3331 329 -3230 330
rect -3331 317 -3330 329
tri -3330 325 -3326 329 ne
tri -3235 325 -3231 329 nw
rect -3231 317 -3230 329
rect -2534 330 -2533 343
tri -2533 330 -2529 334 se
tri -2470 330 -2466 334 sw
rect -2466 330 -2465 343
rect -2534 329 -2465 330
rect -2534 317 -2533 329
tri -2533 325 -2529 329 ne
tri -2470 325 -2466 329 nw
rect -2466 317 -2465 329
rect -2331 330 -2330 343
tri -2330 330 -2326 334 se
tri -2235 330 -2231 334 sw
rect -2231 330 -2230 343
rect -2331 329 -2230 330
rect -2331 317 -2330 329
tri -2330 325 -2326 329 ne
tri -2235 325 -2231 329 nw
rect -2231 317 -2230 329
rect -1534 330 -1533 343
tri -1533 330 -1529 334 se
tri -1470 330 -1466 334 sw
rect -1466 330 -1465 343
rect -1534 329 -1465 330
rect -1534 317 -1533 329
tri -1533 325 -1529 329 ne
tri -1470 325 -1466 329 nw
rect -1466 317 -1465 329
rect -1331 330 -1330 343
tri -1330 330 -1326 334 se
tri -1235 330 -1231 334 sw
rect -1231 330 -1230 343
rect -1331 329 -1230 330
rect -1331 317 -1330 329
tri -1330 325 -1326 329 ne
tri -1235 325 -1231 329 nw
rect -1231 317 -1230 329
rect -534 330 -533 343
tri -533 330 -529 334 se
tri -470 330 -466 334 sw
rect -466 330 -465 343
rect -534 329 -465 330
rect -534 317 -533 329
tri -533 325 -529 329 ne
tri -470 325 -466 329 nw
rect -466 317 -465 329
rect -331 330 -330 343
tri -330 330 -326 334 se
tri -235 330 -231 334 sw
rect -231 330 -230 343
rect -331 329 -230 330
rect -331 317 -330 329
tri -330 325 -326 329 ne
tri -235 325 -231 329 nw
rect -231 317 -230 329
rect 1466 330 1467 343
tri 1467 330 1471 334 se
tri 1530 330 1534 334 sw
rect 1534 330 1535 343
rect 1466 329 1535 330
rect 1466 317 1467 329
tri 1467 325 1471 329 ne
tri 1530 325 1534 329 nw
rect 1534 317 1535 329
rect 1669 330 1670 343
tri 1670 330 1674 334 se
tri 1765 330 1769 334 sw
rect 1769 330 1770 343
rect 1669 329 1770 330
rect 1669 317 1670 329
tri 1670 325 1674 329 ne
tri 1765 325 1769 329 nw
rect 1769 317 1770 329
rect 2466 330 2467 343
tri 2467 330 2471 334 se
tri 2530 330 2534 334 sw
rect 2534 330 2535 343
rect 2466 329 2535 330
rect 2466 317 2467 329
tri 2467 325 2471 329 ne
tri 2530 325 2534 329 nw
rect 2534 317 2535 329
rect 2669 330 2670 343
tri 2670 330 2674 334 se
tri 2765 330 2769 334 sw
rect 2769 330 2770 343
rect 2669 329 2770 330
rect 2669 317 2670 329
tri 2670 325 2674 329 ne
tri 2765 325 2769 329 nw
rect 2769 317 2770 329
rect 3466 330 3467 343
tri 3467 330 3471 334 se
tri 3530 330 3534 334 sw
rect 3534 330 3535 343
rect 3466 329 3535 330
rect 3466 317 3467 329
tri 3467 325 3471 329 ne
tri 3530 325 3534 329 nw
rect 3534 317 3535 329
rect 3669 330 3670 343
tri 3670 330 3674 334 se
tri 3765 330 3769 334 sw
rect 3769 330 3770 343
rect 3669 329 3770 330
rect 3669 317 3670 329
tri 3670 325 3674 329 ne
tri 3765 325 3769 329 nw
rect 3769 317 3770 329
rect -3811 176 -3810 189
tri -3810 176 -3806 180 se
tri -3398 176 -3394 180 sw
rect -3394 176 -3393 189
rect -3811 175 -3623 176
rect -3581 175 -3393 176
rect -3811 163 -3810 175
tri -3810 171 -3806 175 ne
tri -3398 171 -3394 175 nw
rect -3394 163 -3393 175
rect -2811 176 -2810 189
tri -2810 176 -2806 180 se
tri -2398 176 -2394 180 sw
rect -2394 176 -2393 189
rect -2811 175 -2623 176
rect -2581 175 -2393 176
rect -2811 163 -2810 175
tri -2810 171 -2806 175 ne
tri -2398 171 -2394 175 nw
rect -2394 163 -2393 175
rect -1811 176 -1810 189
tri -1810 176 -1806 180 se
tri -1398 176 -1394 180 sw
rect -1394 176 -1393 189
rect -1811 175 -1623 176
rect -1581 175 -1393 176
rect -1811 163 -1810 175
tri -1810 171 -1806 175 ne
tri -1398 171 -1394 175 nw
rect -1394 163 -1393 175
rect -811 176 -810 189
tri -810 176 -806 180 se
tri -398 176 -394 180 sw
rect -394 176 -393 189
rect -811 175 -623 176
rect -581 175 -393 176
rect -811 163 -810 175
tri -810 171 -806 175 ne
tri -398 171 -394 175 nw
rect -394 163 -393 175
rect 1189 176 1190 189
tri 1190 176 1194 180 se
tri 1602 176 1606 180 sw
rect 1606 176 1607 189
rect 1189 175 1377 176
rect 1419 175 1607 176
rect 1189 163 1190 175
tri 1190 171 1194 175 ne
tri 1602 171 1606 175 nw
rect 1606 163 1607 175
rect 2189 176 2190 189
tri 2190 176 2194 180 se
tri 2602 176 2606 180 sw
rect 2606 176 2607 189
rect 2189 175 2377 176
rect 2419 175 2607 176
rect 2189 163 2190 175
tri 2190 171 2194 175 ne
tri 2602 171 2606 175 nw
rect 2606 163 2607 175
rect 3189 176 3190 189
tri 3190 176 3194 180 se
tri 3602 176 3606 180 sw
rect 3606 176 3607 189
rect 3189 175 3377 176
rect 3419 175 3607 176
rect 3189 163 3190 175
tri 3190 171 3194 175 ne
tri 3602 171 3606 175 nw
rect 3606 163 3607 175
rect -3638 136 -3637 149
tri -3637 136 -3633 140 se
tri -3571 136 -3567 140 sw
rect -3567 136 -3566 149
rect -3638 135 -3566 136
rect -3638 123 -3637 135
tri -3637 131 -3633 135 ne
tri -3571 131 -3567 135 nw
rect -3567 123 -3566 135
rect -2638 136 -2637 149
tri -2637 136 -2633 140 se
tri -2571 136 -2567 140 sw
rect -2567 136 -2566 149
rect -2638 135 -2566 136
rect -2638 123 -2637 135
tri -2637 131 -2633 135 ne
tri -2571 131 -2567 135 nw
rect -2567 123 -2566 135
rect -1638 136 -1637 149
tri -1637 136 -1633 140 se
tri -1571 136 -1567 140 sw
rect -1567 136 -1566 149
rect -1638 135 -1566 136
rect -1638 123 -1637 135
tri -1637 131 -1633 135 ne
tri -1571 131 -1567 135 nw
rect -1567 123 -1566 135
rect -638 136 -637 149
tri -637 136 -633 140 se
tri -571 136 -567 140 sw
rect -567 136 -566 149
rect -638 135 -566 136
rect -638 123 -637 135
tri -637 131 -633 135 ne
tri -571 131 -567 135 nw
rect -567 123 -566 135
rect 1362 136 1363 149
tri 1363 136 1367 140 se
tri 1429 136 1433 140 sw
rect 1433 136 1434 149
rect 1362 135 1434 136
rect 1362 123 1363 135
tri 1363 131 1367 135 ne
tri 1429 131 1433 135 nw
rect 1433 123 1434 135
rect 2362 136 2363 149
tri 2363 136 2367 140 se
tri 2429 136 2433 140 sw
rect 2433 136 2434 149
rect 2362 135 2434 136
rect 2362 123 2363 135
tri 2363 131 2367 135 ne
tri 2429 131 2433 135 nw
rect 2433 123 2434 135
rect 3362 136 3363 149
tri 3363 136 3367 140 se
tri 3429 136 3433 140 sw
rect 3433 136 3434 149
rect 3362 135 3434 136
rect 3362 123 3363 135
tri 3363 131 3367 135 ne
tri 3429 131 3433 135 nw
rect 3433 123 3434 135
rect -3974 -217 -3973 -204
tri -3973 -217 -3969 -213 se
tri -3235 -217 -3231 -213 sw
rect -3231 -217 -3230 -204
rect -3974 -218 -3629 -217
rect -3576 -218 -3230 -217
rect -3974 -230 -3973 -218
tri -3973 -222 -3969 -218 ne
tri -3235 -222 -3231 -218 nw
rect -3231 -230 -3230 -218
rect -2974 -217 -2973 -204
tri -2973 -217 -2969 -213 se
tri -2235 -217 -2231 -213 sw
rect -2231 -217 -2230 -204
rect -2974 -218 -2629 -217
rect -2576 -218 -2230 -217
rect -2974 -230 -2973 -218
tri -2973 -222 -2969 -218 ne
tri -2235 -222 -2231 -218 nw
rect -2231 -230 -2230 -218
rect -1974 -217 -1973 -204
tri -1973 -217 -1969 -213 se
tri -1235 -217 -1231 -213 sw
rect -1231 -217 -1230 -204
rect -1974 -218 -1629 -217
rect -1576 -218 -1230 -217
rect -1974 -230 -1973 -218
tri -1973 -222 -1969 -218 ne
tri -1235 -222 -1231 -218 nw
rect -1231 -230 -1230 -218
rect -974 -217 -973 -204
tri -973 -217 -969 -213 se
tri -235 -217 -231 -213 sw
rect -231 -217 -230 -204
rect -974 -218 -629 -217
rect -576 -218 -230 -217
rect -974 -230 -973 -218
tri -973 -222 -969 -218 ne
tri -235 -222 -231 -218 nw
rect -231 -230 -230 -218
rect 26 -217 27 -204
tri 27 -217 31 -213 se
tri 765 -217 769 -213 sw
rect 769 -217 770 -204
rect 26 -218 371 -217
rect 424 -218 770 -217
rect 26 -230 27 -218
tri 27 -222 31 -218 ne
tri 765 -222 769 -218 nw
rect 769 -230 770 -218
rect 1026 -217 1027 -204
tri 1027 -217 1031 -213 se
tri 1765 -217 1769 -213 sw
rect 1769 -217 1770 -204
rect 1026 -218 1371 -217
rect 1424 -218 1770 -217
rect 1026 -230 1027 -218
tri 1027 -222 1031 -218 ne
tri 1765 -222 1769 -218 nw
rect 1769 -230 1770 -218
rect 2026 -217 2027 -204
tri 2027 -217 2031 -213 se
tri 2765 -217 2769 -213 sw
rect 2769 -217 2770 -204
rect 2026 -218 2371 -217
rect 2424 -218 2770 -217
rect 2026 -230 2027 -218
tri 2027 -222 2031 -218 ne
tri 2765 -222 2769 -218 nw
rect 2769 -230 2770 -218
rect 3026 -217 3027 -204
tri 3027 -217 3031 -213 se
tri 3765 -217 3769 -213 sw
rect 3769 -217 3770 -204
rect 3026 -218 3371 -217
rect 3424 -218 3770 -217
rect 3026 -230 3027 -218
tri 3027 -222 3031 -218 ne
tri 3765 -222 3769 -218 nw
rect 3769 -230 3770 -218
rect -3847 -380 -3846 -367
tri -3846 -380 -3842 -376 se
tri -3362 -380 -3358 -376 sw
rect -3358 -380 -3357 -367
rect -3847 -381 -3655 -380
rect -3548 -381 -3357 -380
rect -3847 -393 -3846 -381
tri -3846 -385 -3842 -381 ne
tri -3362 -385 -3358 -381 nw
rect -3358 -393 -3357 -381
rect -2847 -380 -2846 -367
tri -2846 -380 -2842 -376 se
tri -2362 -380 -2358 -376 sw
rect -2358 -380 -2357 -367
rect -2847 -381 -2655 -380
rect -2548 -381 -2357 -380
rect -2847 -393 -2846 -381
tri -2846 -385 -2842 -381 ne
tri -2362 -385 -2358 -381 nw
rect -2358 -393 -2357 -381
rect -1847 -380 -1846 -367
tri -1846 -380 -1842 -376 se
tri -1362 -380 -1358 -376 sw
rect -1358 -380 -1357 -367
rect -1847 -381 -1655 -380
rect -1548 -381 -1357 -380
rect -1847 -393 -1846 -381
tri -1846 -385 -1842 -381 ne
tri -1362 -385 -1358 -381 nw
rect -1358 -393 -1357 -381
rect -847 -380 -846 -367
tri -846 -380 -842 -376 se
tri -362 -380 -358 -376 sw
rect -358 -380 -357 -367
rect -847 -381 -655 -380
rect -548 -381 -357 -380
rect -847 -393 -846 -381
tri -846 -385 -842 -381 ne
tri -362 -385 -358 -381 nw
rect -358 -393 -357 -381
rect 153 -380 154 -367
tri 154 -380 158 -376 se
tri 638 -380 642 -376 sw
rect 642 -380 643 -367
rect 153 -381 345 -380
rect 452 -381 643 -380
rect 153 -393 154 -381
tri 154 -385 158 -381 ne
tri 638 -385 642 -381 nw
rect 642 -393 643 -381
rect 1153 -380 1154 -367
tri 1154 -380 1158 -376 se
tri 1638 -380 1642 -376 sw
rect 1642 -380 1643 -367
rect 1153 -381 1345 -380
rect 1452 -381 1643 -380
rect 1153 -393 1154 -381
tri 1154 -385 1158 -381 ne
tri 1638 -385 1642 -381 nw
rect 1642 -393 1643 -381
rect 2153 -380 2154 -367
tri 2154 -380 2158 -376 se
tri 2638 -380 2642 -376 sw
rect 2642 -380 2643 -367
rect 2153 -381 2345 -380
rect 2452 -381 2643 -380
rect 2153 -393 2154 -381
tri 2154 -385 2158 -381 ne
tri 2638 -385 2642 -381 nw
rect 2642 -393 2643 -381
rect 3153 -380 3154 -367
tri 3154 -380 3158 -376 se
tri 3638 -380 3642 -376 sw
rect 3642 -380 3643 -367
rect 3153 -381 3345 -380
rect 3452 -381 3643 -380
rect 3153 -393 3154 -381
tri 3154 -385 3158 -381 ne
tri 3638 -385 3642 -381 nw
rect 3642 -393 3643 -381
rect -3811 -435 -3810 -422
tri -3810 -435 -3806 -431 se
tri -3792 -435 -3788 -431 sw
rect -3788 -435 -3787 -422
rect -3811 -436 -3787 -435
rect -3811 -448 -3810 -436
tri -3810 -440 -3806 -436 ne
tri -3801 -440 -3799 -437 se
tri -3792 -440 -3788 -436 nw
tri -3802 -443 -3801 -440 se
rect -3801 -443 -3799 -440
tri -3799 -443 -3798 -440 sw
rect -3803 -444 -3802 -443
tri -3802 -444 -3801 -443 nw
rect -3799 -444 -3798 -443
rect -3805 -476 -3800 -444
rect -3788 -448 -3787 -436
rect -2811 -435 -2810 -422
tri -2810 -435 -2806 -431 se
tri -2792 -435 -2788 -431 sw
rect -2788 -435 -2787 -422
rect -2811 -436 -2787 -435
rect -2811 -448 -2810 -436
tri -2810 -440 -2806 -436 ne
tri -2801 -440 -2799 -437 se
tri -2802 -443 -2801 -440 se
rect -2801 -443 -2799 -440
tri -2799 -443 -2798 -437 sw
tri -2792 -440 -2788 -436 nw
rect -2803 -444 -2802 -443
tri -2802 -444 -2801 -443 nw
rect -2799 -444 -2798 -443
rect -3393 -467 -3392 -454
tri -3392 -467 -3388 -463 se
tri -3336 -467 -3332 -463 sw
rect -3332 -467 -3331 -454
rect -3393 -468 -3331 -467
rect -3393 -480 -3392 -468
tri -3392 -472 -3388 -468 ne
tri -3336 -472 -3332 -468 nw
rect -3332 -480 -3331 -468
rect -2805 -476 -2800 -444
rect -2788 -448 -2787 -436
rect -1811 -435 -1810 -422
tri -1810 -435 -1806 -431 se
tri -1792 -435 -1788 -431 sw
rect -1788 -435 -1787 -422
rect -1811 -436 -1787 -435
rect -1811 -448 -1810 -436
tri -1810 -440 -1806 -436 ne
tri -1801 -440 -1799 -437 se
tri -1792 -440 -1788 -436 nw
tri -1802 -443 -1801 -440 se
rect -1801 -443 -1799 -440
tri -1799 -443 -1798 -440 sw
rect -1803 -444 -1802 -443
tri -1802 -444 -1801 -443 nw
rect -1799 -444 -1798 -443
rect -2393 -467 -2392 -454
tri -2392 -467 -2388 -463 se
tri -2336 -467 -2332 -463 sw
rect -2332 -467 -2331 -454
rect -2393 -468 -2331 -467
rect -2393 -480 -2392 -468
tri -2392 -472 -2388 -468 ne
tri -2336 -472 -2332 -468 nw
rect -2332 -480 -2331 -468
rect -1805 -476 -1800 -444
rect -1788 -448 -1787 -436
rect -811 -435 -810 -422
tri -810 -435 -806 -431 se
tri -792 -435 -788 -431 sw
rect -788 -435 -787 -422
rect -811 -436 -787 -435
rect -811 -448 -810 -436
tri -810 -440 -806 -436 ne
tri -801 -440 -799 -437 se
tri -792 -440 -788 -436 nw
tri -802 -443 -801 -440 se
rect -801 -443 -799 -440
tri -799 -443 -798 -440 sw
rect -803 -444 -802 -443
tri -802 -444 -801 -443 nw
rect -799 -444 -798 -443
rect -1393 -467 -1392 -454
tri -1392 -467 -1388 -463 se
tri -1336 -467 -1332 -463 sw
rect -1332 -467 -1331 -454
rect -1393 -468 -1331 -467
rect -1393 -480 -1392 -468
tri -1392 -472 -1388 -468 ne
tri -1336 -472 -1332 -468 nw
rect -1332 -480 -1331 -468
rect -805 -476 -800 -444
rect -788 -448 -787 -436
rect 189 -435 190 -422
tri 190 -435 194 -431 se
tri 208 -435 212 -431 sw
rect 212 -435 213 -422
rect 189 -436 213 -435
rect 189 -448 190 -436
tri 190 -440 194 -436 ne
tri 199 -440 201 -437 se
tri 198 -443 199 -440 se
rect 199 -443 201 -440
tri 201 -443 202 -437 sw
tri 208 -440 212 -436 nw
rect 197 -444 198 -443
tri 198 -444 199 -443 nw
rect 201 -444 202 -443
rect -393 -467 -392 -454
tri -392 -467 -388 -463 se
tri -336 -467 -332 -463 sw
rect -332 -467 -331 -454
rect -393 -468 -331 -467
rect -393 -480 -392 -468
tri -392 -472 -388 -468 ne
tri -336 -472 -332 -468 nw
rect -332 -480 -331 -468
rect 195 -476 200 -444
rect 212 -448 213 -436
rect 1189 -435 1190 -422
tri 1190 -435 1194 -431 se
tri 1208 -435 1212 -431 sw
rect 1212 -435 1213 -422
rect 1189 -436 1213 -435
rect 1189 -448 1190 -436
tri 1190 -440 1194 -436 ne
tri 1199 -440 1201 -437 se
tri 1208 -440 1212 -436 nw
tri 1198 -443 1199 -440 se
rect 1199 -443 1201 -440
tri 1201 -443 1202 -440 sw
rect 1197 -444 1198 -443
tri 1198 -444 1199 -443 nw
rect 1201 -444 1202 -443
rect 607 -467 608 -454
tri 608 -467 612 -463 se
tri 664 -467 668 -463 sw
rect 668 -467 669 -454
rect 607 -468 669 -467
rect 607 -480 608 -468
tri 608 -472 612 -468 ne
tri 664 -472 668 -468 nw
rect 668 -480 669 -468
rect 1195 -476 1200 -444
rect 1212 -448 1213 -436
rect 2189 -435 2190 -422
tri 2190 -435 2194 -431 se
tri 2208 -435 2212 -431 sw
rect 2212 -435 2213 -422
rect 2189 -436 2213 -435
rect 2189 -448 2190 -436
tri 2190 -440 2194 -436 ne
tri 2199 -440 2201 -437 se
tri 2208 -440 2212 -436 nw
tri 2198 -443 2199 -440 se
rect 2199 -443 2201 -440
tri 2201 -443 2202 -440 sw
rect 2197 -444 2198 -443
tri 2198 -444 2199 -443 nw
rect 2201 -444 2202 -443
rect 1607 -467 1608 -454
tri 1608 -467 1612 -463 se
tri 1664 -467 1668 -463 sw
rect 1668 -467 1669 -454
rect 1607 -468 1669 -467
rect 1607 -480 1608 -468
tri 1608 -472 1612 -468 ne
tri 1664 -472 1668 -468 nw
rect 1668 -480 1669 -468
rect 2195 -476 2200 -444
rect 2212 -448 2213 -436
rect 3189 -435 3190 -422
tri 3190 -435 3194 -431 se
tri 3208 -435 3212 -431 sw
rect 3212 -435 3213 -422
rect 3189 -436 3213 -435
rect 3189 -448 3190 -436
tri 3190 -440 3194 -436 ne
tri 3199 -440 3201 -437 se
tri 3208 -440 3212 -436 nw
tri 3198 -443 3199 -440 se
rect 3199 -443 3201 -440
tri 3201 -443 3202 -440 sw
rect 3197 -444 3198 -443
tri 3198 -444 3199 -443 nw
rect 3201 -444 3202 -443
rect 2607 -467 2608 -454
tri 2608 -467 2612 -463 se
tri 2664 -467 2668 -463 sw
rect 2668 -467 2669 -454
rect 2607 -468 2669 -467
rect 2607 -480 2608 -468
tri 2608 -472 2612 -468 ne
tri 2664 -472 2668 -468 nw
rect 2668 -480 2669 -468
rect 3195 -476 3200 -444
rect 3212 -448 3213 -436
rect 3607 -467 3608 -454
tri 3608 -467 3612 -463 se
tri 3664 -467 3668 -463 sw
rect 3668 -467 3669 -454
rect 3607 -468 3669 -467
rect 3607 -480 3608 -468
tri 3608 -472 3612 -468 ne
tri 3664 -472 3668 -468 nw
rect 3668 -480 3669 -468
rect -3670 -521 -3669 -508
tri -3669 -521 -3665 -517 se
tri -3539 -521 -3535 -517 sw
rect -3535 -521 -3534 -508
rect -3670 -522 -3623 -521
rect -3581 -522 -3534 -521
rect -3670 -534 -3669 -522
tri -3669 -526 -3665 -522 ne
tri -3539 -526 -3535 -522 nw
rect -3535 -534 -3534 -522
rect -2670 -521 -2669 -508
tri -2669 -521 -2665 -517 se
tri -2539 -521 -2535 -517 sw
rect -2535 -521 -2534 -508
rect -2670 -522 -2623 -521
rect -2581 -522 -2534 -521
rect -2670 -534 -2669 -522
tri -2669 -526 -2665 -522 ne
tri -2539 -526 -2535 -522 nw
rect -2535 -534 -2534 -522
rect -1670 -521 -1669 -508
tri -1669 -521 -1665 -517 se
tri -1539 -521 -1535 -517 sw
rect -1535 -521 -1534 -508
rect -1670 -522 -1623 -521
rect -1581 -522 -1534 -521
rect -1670 -534 -1669 -522
tri -1669 -526 -1665 -522 ne
tri -1539 -526 -1535 -522 nw
rect -1535 -534 -1534 -522
rect -670 -521 -669 -508
tri -669 -521 -665 -517 se
tri -539 -521 -535 -517 sw
rect -535 -521 -534 -508
rect -670 -522 -623 -521
rect -581 -522 -534 -521
rect -670 -534 -669 -522
tri -669 -526 -665 -522 ne
tri -539 -526 -535 -522 nw
rect -535 -534 -534 -522
rect 330 -521 331 -508
tri 331 -521 335 -517 se
tri 461 -521 465 -517 sw
rect 465 -521 466 -508
rect 330 -522 377 -521
rect 419 -522 466 -521
rect 330 -534 331 -522
tri 331 -526 335 -522 ne
tri 461 -526 465 -522 nw
rect 465 -534 466 -522
rect 1330 -521 1331 -508
tri 1331 -521 1335 -517 se
tri 1461 -521 1465 -517 sw
rect 1465 -521 1466 -508
rect 1330 -522 1377 -521
rect 1419 -522 1466 -521
rect 1330 -534 1331 -522
tri 1331 -526 1335 -522 ne
tri 1461 -526 1465 -522 nw
rect 1465 -534 1466 -522
rect 2330 -521 2331 -508
tri 2331 -521 2335 -517 se
tri 2461 -521 2465 -517 sw
rect 2465 -521 2466 -508
rect 2330 -522 2377 -521
rect 2419 -522 2466 -521
rect 2330 -534 2331 -522
tri 2331 -526 2335 -522 ne
tri 2461 -526 2465 -522 nw
rect 2465 -534 2466 -522
rect 3330 -521 3331 -508
tri 3331 -521 3335 -517 se
tri 3461 -521 3465 -517 sw
rect 3465 -521 3466 -508
rect 3330 -522 3377 -521
rect 3419 -522 3466 -521
rect 3330 -534 3331 -522
tri 3331 -526 3335 -522 ne
tri 3461 -526 3465 -522 nw
rect 3465 -534 3466 -522
rect -3811 -558 -3810 -545
tri -3810 -558 -3806 -554 se
tri -3744 -558 -3740 -554 sw
rect -3740 -558 -3739 -545
rect -3811 -559 -3739 -558
rect -3811 -571 -3810 -559
tri -3810 -563 -3806 -559 ne
tri -3744 -563 -3740 -559 nw
rect -3740 -571 -3739 -559
rect -2811 -558 -2810 -545
tri -2810 -558 -2806 -554 se
tri -2744 -558 -2740 -554 sw
rect -2740 -558 -2739 -545
rect -2811 -559 -2739 -558
rect -2811 -571 -2810 -559
tri -2810 -563 -2806 -559 ne
tri -2744 -563 -2740 -559 nw
rect -2740 -571 -2739 -559
rect -1811 -558 -1810 -545
tri -1810 -558 -1806 -554 se
tri -1744 -558 -1740 -554 sw
rect -1740 -558 -1739 -545
rect -1811 -559 -1739 -558
rect -1811 -571 -1810 -559
tri -1810 -563 -1806 -559 ne
tri -1744 -563 -1740 -559 nw
rect -1740 -571 -1739 -559
rect -811 -558 -810 -545
tri -810 -558 -806 -554 se
tri -744 -558 -740 -554 sw
rect -740 -558 -739 -545
rect -811 -559 -739 -558
rect -811 -571 -810 -559
tri -810 -563 -806 -559 ne
tri -744 -563 -740 -559 nw
rect -740 -571 -739 -559
rect 189 -558 190 -545
tri 190 -558 194 -554 se
tri 256 -558 260 -554 sw
rect 260 -558 261 -545
rect 189 -559 261 -558
rect 189 -571 190 -559
tri 190 -563 194 -559 ne
tri 256 -563 260 -559 nw
rect 260 -571 261 -559
rect 1189 -558 1190 -545
tri 1190 -558 1194 -554 se
tri 1256 -558 1260 -554 sw
rect 1260 -558 1261 -545
rect 1189 -559 1261 -558
rect 1189 -571 1190 -559
tri 1190 -563 1194 -559 ne
tri 1256 -563 1260 -559 nw
rect 1260 -571 1261 -559
rect 2189 -558 2190 -545
tri 2190 -558 2194 -554 se
tri 2256 -558 2260 -554 sw
rect 2260 -558 2261 -545
rect 2189 -559 2261 -558
rect 2189 -571 2190 -559
tri 2190 -563 2194 -559 ne
tri 2256 -563 2260 -559 nw
rect 2260 -571 2261 -559
rect 3189 -558 3190 -545
tri 3190 -558 3194 -554 se
tri 3256 -558 3260 -554 sw
rect 3260 -558 3261 -545
rect 3189 -559 3261 -558
rect 3189 -571 3190 -559
tri 3190 -563 3194 -559 ne
tri 3256 -563 3260 -559 nw
rect 3260 -571 3261 -559
tri -3610 -596 -3608 -594 se
tri -3608 -596 -3607 -594 sw
tri -3597 -596 -3596 -594 se
tri -3596 -596 -3594 -594 sw
tri -3610 -597 -3608 -596 ne
rect -3608 -597 -3607 -596
tri -3607 -597 -3605 -596 sw
tri -3599 -597 -3597 -596 se
tri -3608 -600 -3605 -597 ne
tri -3605 -599 -3604 -597 sw
tri -3600 -599 -3599 -597 se
rect -3599 -599 -3597 -597
tri -3597 -599 -3594 -596 nw
tri -2610 -596 -2608 -594 se
tri -2608 -596 -2607 -594 sw
tri -2597 -596 -2596 -594 se
tri -2596 -596 -2594 -594 sw
tri -2610 -597 -2608 -596 ne
rect -2608 -597 -2607 -596
tri -2607 -597 -2605 -596 sw
tri -2599 -597 -2597 -596 se
rect -3605 -600 -3604 -599
tri -3604 -600 -3602 -599 sw
tri -3602 -600 -3600 -599 se
tri -3605 -602 -3604 -600 ne
tri -3607 -605 -3604 -602 se
rect -3604 -604 -3600 -600
tri -3600 -602 -3597 -599 nw
tri -2608 -600 -2605 -597 ne
tri -2605 -599 -2604 -597 sw
tri -2600 -599 -2599 -597 se
rect -2599 -599 -2597 -597
tri -2597 -599 -2594 -596 nw
tri -1610 -596 -1608 -594 se
tri -1608 -596 -1607 -594 sw
tri -1597 -596 -1596 -594 se
tri -1596 -596 -1594 -594 sw
tri -1610 -597 -1608 -596 ne
rect -1608 -597 -1607 -596
tri -1607 -597 -1605 -596 sw
tri -1599 -597 -1597 -596 se
rect -2605 -600 -2604 -599
tri -2604 -600 -2602 -599 sw
tri -2602 -600 -2600 -599 se
tri -2605 -602 -2604 -600 ne
rect -3604 -605 -3603 -604
tri -3603 -605 -3602 -604 nw
tri -3602 -605 -3601 -604 ne
rect -3601 -605 -3600 -604
tri -3600 -605 -3597 -602 sw
tri -2607 -605 -2604 -602 se
rect -2604 -604 -2600 -600
tri -2600 -602 -2597 -599 nw
tri -1608 -600 -1605 -597 ne
tri -1605 -599 -1604 -597 sw
tri -1600 -599 -1599 -597 se
rect -1599 -599 -1597 -597
tri -1597 -599 -1594 -596 nw
tri -610 -596 -608 -594 se
tri -608 -596 -607 -594 sw
tri -597 -596 -596 -594 se
tri -596 -596 -594 -594 sw
tri -610 -597 -608 -596 ne
rect -608 -597 -607 -596
tri -607 -597 -605 -596 sw
tri -599 -597 -597 -596 se
rect -1605 -600 -1604 -599
tri -1604 -600 -1602 -599 sw
tri -1602 -600 -1600 -599 se
tri -1605 -602 -1604 -600 ne
rect -2604 -605 -2603 -604
tri -2603 -605 -2602 -604 nw
tri -2602 -605 -2601 -604 ne
rect -2601 -605 -2600 -604
tri -2600 -605 -2597 -602 sw
tri -1607 -605 -1604 -602 se
rect -1604 -604 -1600 -600
tri -1600 -602 -1597 -599 nw
tri -608 -600 -605 -597 ne
tri -605 -599 -604 -597 sw
tri -600 -599 -599 -597 se
rect -599 -599 -597 -597
tri -597 -599 -594 -596 nw
tri 390 -596 392 -594 se
tri 392 -596 393 -594 sw
tri 403 -596 404 -594 se
tri 404 -596 406 -594 sw
tri 390 -597 392 -596 ne
rect 392 -597 393 -596
tri 393 -597 395 -596 sw
tri 401 -597 403 -596 se
rect -605 -600 -604 -599
tri -604 -600 -602 -599 sw
tri -602 -600 -600 -599 se
tri -605 -602 -604 -600 ne
rect -1604 -605 -1603 -604
tri -1603 -605 -1602 -604 nw
tri -1602 -605 -1601 -604 ne
rect -1601 -605 -1600 -604
tri -1600 -605 -1597 -602 sw
tri -607 -605 -604 -602 se
rect -604 -604 -600 -600
tri -600 -602 -597 -599 nw
tri 392 -600 395 -597 ne
tri 395 -599 396 -597 sw
tri 400 -599 401 -597 se
rect 401 -599 403 -597
tri 403 -599 406 -596 nw
tri 1390 -596 1392 -594 se
tri 1392 -596 1393 -594 sw
tri 1403 -596 1404 -594 se
tri 1404 -596 1406 -594 sw
tri 1390 -597 1392 -596 ne
rect 1392 -597 1393 -596
tri 1393 -597 1395 -596 sw
tri 1401 -597 1403 -596 se
rect 395 -600 396 -599
tri 396 -600 398 -599 sw
tri 398 -600 400 -599 se
tri 395 -602 396 -600 ne
rect -604 -605 -603 -604
tri -603 -605 -602 -604 nw
tri -602 -605 -601 -604 ne
rect -601 -605 -600 -604
tri -600 -605 -597 -602 sw
tri 393 -605 396 -602 se
rect 396 -604 400 -600
tri 400 -602 403 -599 nw
tri 1392 -600 1395 -597 ne
tri 1395 -599 1396 -597 sw
tri 1400 -599 1401 -597 se
rect 1401 -599 1403 -597
tri 1403 -599 1406 -596 nw
tri 2390 -596 2392 -594 se
tri 2392 -596 2393 -594 sw
tri 2403 -596 2404 -594 se
tri 2404 -596 2406 -594 sw
tri 2390 -597 2392 -596 ne
rect 2392 -597 2393 -596
tri 2393 -597 2395 -596 sw
tri 2401 -597 2403 -596 se
rect 1395 -600 1396 -599
tri 1396 -600 1398 -599 sw
tri 1398 -600 1400 -599 se
tri 1395 -602 1396 -600 ne
rect 396 -605 397 -604
tri 397 -605 398 -604 nw
tri 398 -605 399 -604 ne
rect 399 -605 400 -604
tri 400 -605 403 -602 sw
tri 1393 -605 1396 -602 se
rect 1396 -604 1400 -600
tri 1400 -602 1403 -599 nw
tri 2392 -600 2395 -597 ne
tri 2395 -599 2396 -597 sw
tri 2400 -599 2401 -597 se
rect 2401 -599 2403 -597
tri 2403 -599 2406 -596 nw
tri 3390 -596 3392 -594 se
tri 3392 -596 3393 -594 sw
tri 3403 -596 3404 -594 se
tri 3404 -596 3406 -594 sw
tri 3390 -597 3392 -596 ne
rect 3392 -597 3393 -596
tri 3393 -597 3395 -596 sw
tri 3401 -597 3403 -596 se
rect 2395 -600 2396 -599
tri 2396 -600 2398 -599 sw
tri 2398 -600 2400 -599 se
tri 2395 -602 2396 -600 ne
rect 1396 -605 1397 -604
tri 1397 -605 1398 -604 nw
tri 1398 -605 1399 -604 ne
rect 1399 -605 1400 -604
tri 1400 -605 1403 -602 sw
tri 2393 -605 2396 -602 se
rect 2396 -604 2400 -600
tri 2400 -602 2403 -599 nw
tri 3392 -600 3395 -597 ne
tri 3395 -599 3396 -597 sw
tri 3400 -599 3401 -597 se
rect 3401 -599 3403 -597
tri 3403 -599 3406 -596 nw
rect 3395 -600 3396 -599
tri 3396 -600 3398 -599 sw
tri 3398 -600 3400 -599 se
tri 3395 -602 3396 -600 ne
rect 2396 -605 2397 -604
tri 2397 -605 2398 -604 nw
tri 2398 -605 2399 -604 ne
rect 2399 -605 2400 -604
tri 2400 -605 2403 -602 sw
tri 3393 -605 3396 -602 se
rect 3396 -604 3400 -600
tri 3400 -602 3403 -599 nw
rect 3396 -605 3397 -604
tri 3397 -605 3398 -604 nw
tri 3398 -605 3399 -604 ne
rect 3399 -605 3400 -604
tri 3400 -605 3403 -602 sw
tri -3610 -608 -3607 -605 se
tri -3607 -608 -3604 -605 nw
tri -3600 -608 -3597 -605 ne
tri -3597 -608 -3594 -605 sw
tri -3610 -610 -3608 -608 ne
tri -3608 -610 -3607 -608 nw
tri -3597 -610 -3596 -608 ne
tri -3596 -610 -3594 -608 nw
tri -2610 -608 -2607 -605 se
tri -2607 -608 -2604 -605 nw
tri -2600 -608 -2597 -605 ne
tri -2597 -608 -2594 -605 sw
tri -2610 -610 -2608 -608 ne
tri -2608 -610 -2607 -608 nw
tri -2597 -610 -2596 -608 ne
tri -2596 -610 -2594 -608 nw
tri -1610 -608 -1607 -605 se
tri -1607 -608 -1604 -605 nw
tri -1600 -608 -1597 -605 ne
tri -1597 -608 -1594 -605 sw
tri -1610 -610 -1608 -608 ne
tri -1608 -610 -1607 -608 nw
tri -1597 -610 -1596 -608 ne
tri -1596 -610 -1594 -608 nw
tri -610 -608 -607 -605 se
tri -607 -608 -604 -605 nw
tri -600 -608 -597 -605 ne
tri -597 -608 -594 -605 sw
tri -610 -610 -608 -608 ne
tri -608 -610 -607 -608 nw
tri -597 -610 -596 -608 ne
tri -596 -610 -594 -608 nw
tri 390 -608 393 -605 se
tri 393 -608 396 -605 nw
tri 400 -608 403 -605 ne
tri 403 -608 406 -605 sw
tri 390 -610 392 -608 ne
tri 392 -610 393 -608 nw
tri 403 -610 404 -608 ne
tri 404 -610 406 -608 nw
tri 1390 -608 1393 -605 se
tri 1393 -608 1396 -605 nw
tri 1400 -608 1403 -605 ne
tri 1403 -608 1406 -605 sw
tri 1390 -610 1392 -608 ne
tri 1392 -610 1393 -608 nw
tri 1403 -610 1404 -608 ne
tri 1404 -610 1406 -608 nw
tri 2390 -608 2393 -605 se
tri 2393 -608 2396 -605 nw
tri 2400 -608 2403 -605 ne
tri 2403 -608 2406 -605 sw
tri 2390 -610 2392 -608 ne
tri 2392 -610 2393 -608 nw
tri 2403 -610 2404 -608 ne
tri 2404 -610 2406 -608 nw
tri 3390 -608 3393 -605 se
tri 3393 -608 3396 -605 nw
tri 3400 -608 3403 -605 ne
tri 3403 -608 3406 -605 sw
tri 3390 -610 3392 -608 ne
tri 3392 -610 3393 -608 nw
tri 3403 -610 3404 -608 ne
tri 3404 -610 3406 -608 nw
rect -3534 -670 -3533 -657
tri -3533 -670 -3529 -666 se
tri -3470 -670 -3466 -666 sw
rect -3466 -670 -3465 -657
rect -3534 -671 -3465 -670
rect -3534 -683 -3533 -671
tri -3533 -675 -3529 -671 ne
tri -3470 -675 -3466 -671 nw
rect -3466 -683 -3465 -671
rect -3331 -670 -3330 -657
tri -3330 -670 -3326 -666 se
tri -3235 -670 -3231 -666 sw
rect -3231 -670 -3230 -657
rect -3331 -671 -3230 -670
rect -3331 -683 -3330 -671
tri -3330 -675 -3326 -671 ne
tri -3235 -675 -3231 -671 nw
rect -3231 -683 -3230 -671
rect -2534 -670 -2533 -657
tri -2533 -670 -2529 -666 se
tri -2470 -670 -2466 -666 sw
rect -2466 -670 -2465 -657
rect -2534 -671 -2465 -670
rect -2534 -683 -2533 -671
tri -2533 -675 -2529 -671 ne
tri -2470 -675 -2466 -671 nw
rect -2466 -683 -2465 -671
rect -2331 -670 -2330 -657
tri -2330 -670 -2326 -666 se
tri -2235 -670 -2231 -666 sw
rect -2231 -670 -2230 -657
rect -2331 -671 -2230 -670
rect -2331 -683 -2330 -671
tri -2330 -675 -2326 -671 ne
tri -2235 -675 -2231 -671 nw
rect -2231 -683 -2230 -671
rect -1534 -670 -1533 -657
tri -1533 -670 -1529 -666 se
tri -1470 -670 -1466 -666 sw
rect -1466 -670 -1465 -657
rect -1534 -671 -1465 -670
rect -1534 -683 -1533 -671
tri -1533 -675 -1529 -671 ne
tri -1470 -675 -1466 -671 nw
rect -1466 -683 -1465 -671
rect -1331 -670 -1330 -657
tri -1330 -670 -1326 -666 se
tri -1235 -670 -1231 -666 sw
rect -1231 -670 -1230 -657
rect -1331 -671 -1230 -670
rect -1331 -683 -1330 -671
tri -1330 -675 -1326 -671 ne
tri -1235 -675 -1231 -671 nw
rect -1231 -683 -1230 -671
rect -534 -670 -533 -657
tri -533 -670 -529 -666 se
tri -470 -670 -466 -666 sw
rect -466 -670 -465 -657
rect -534 -671 -465 -670
rect -534 -683 -533 -671
tri -533 -675 -529 -671 ne
tri -470 -675 -466 -671 nw
rect -466 -683 -465 -671
rect -331 -670 -330 -657
tri -330 -670 -326 -666 se
tri -235 -670 -231 -666 sw
rect -231 -670 -230 -657
rect -331 -671 -230 -670
rect -331 -683 -330 -671
tri -330 -675 -326 -671 ne
tri -235 -675 -231 -671 nw
rect -231 -683 -230 -671
rect 466 -670 467 -657
tri 467 -670 471 -666 se
tri 530 -670 534 -666 sw
rect 534 -670 535 -657
rect 466 -671 535 -670
rect 466 -683 467 -671
tri 467 -675 471 -671 ne
tri 530 -675 534 -671 nw
rect 534 -683 535 -671
rect 669 -670 670 -657
tri 670 -670 674 -666 se
tri 765 -670 769 -666 sw
rect 769 -670 770 -657
rect 669 -671 770 -670
rect 669 -683 670 -671
tri 670 -675 674 -671 ne
tri 765 -675 769 -671 nw
rect 769 -683 770 -671
rect 1466 -670 1467 -657
tri 1467 -670 1471 -666 se
tri 1530 -670 1534 -666 sw
rect 1534 -670 1535 -657
rect 1466 -671 1535 -670
rect 1466 -683 1467 -671
tri 1467 -675 1471 -671 ne
tri 1530 -675 1534 -671 nw
rect 1534 -683 1535 -671
rect 1669 -670 1670 -657
tri 1670 -670 1674 -666 se
tri 1765 -670 1769 -666 sw
rect 1769 -670 1770 -657
rect 1669 -671 1770 -670
rect 1669 -683 1670 -671
tri 1670 -675 1674 -671 ne
tri 1765 -675 1769 -671 nw
rect 1769 -683 1770 -671
rect 2466 -670 2467 -657
tri 2467 -670 2471 -666 se
tri 2530 -670 2534 -666 sw
rect 2534 -670 2535 -657
rect 2466 -671 2535 -670
rect 2466 -683 2467 -671
tri 2467 -675 2471 -671 ne
tri 2530 -675 2534 -671 nw
rect 2534 -683 2535 -671
rect 2669 -670 2670 -657
tri 2670 -670 2674 -666 se
tri 2765 -670 2769 -666 sw
rect 2769 -670 2770 -657
rect 2669 -671 2770 -670
rect 2669 -683 2670 -671
tri 2670 -675 2674 -671 ne
tri 2765 -675 2769 -671 nw
rect 2769 -683 2770 -671
rect 3466 -670 3467 -657
tri 3467 -670 3471 -666 se
tri 3530 -670 3534 -666 sw
rect 3534 -670 3535 -657
rect 3466 -671 3535 -670
rect 3466 -683 3467 -671
tri 3467 -675 3471 -671 ne
tri 3530 -675 3534 -671 nw
rect 3534 -683 3535 -671
rect 3669 -670 3670 -657
tri 3670 -670 3674 -666 se
tri 3765 -670 3769 -666 sw
rect 3769 -670 3770 -657
rect 3669 -671 3770 -670
rect 3669 -683 3670 -671
tri 3670 -675 3674 -671 ne
tri 3765 -675 3769 -671 nw
rect 3769 -683 3770 -671
rect -3811 -824 -3810 -811
tri -3810 -824 -3806 -820 se
tri -3398 -824 -3394 -820 sw
rect -3394 -824 -3393 -811
rect -3811 -825 -3623 -824
rect -3581 -825 -3393 -824
rect -3811 -837 -3810 -825
tri -3810 -829 -3806 -825 ne
tri -3398 -829 -3394 -825 nw
rect -3394 -837 -3393 -825
rect -2811 -824 -2810 -811
tri -2810 -824 -2806 -820 se
tri -2398 -824 -2394 -820 sw
rect -2394 -824 -2393 -811
rect -2811 -825 -2623 -824
rect -2581 -825 -2393 -824
rect -2811 -837 -2810 -825
tri -2810 -829 -2806 -825 ne
tri -2398 -829 -2394 -825 nw
rect -2394 -837 -2393 -825
rect -1811 -824 -1810 -811
tri -1810 -824 -1806 -820 se
tri -1398 -824 -1394 -820 sw
rect -1394 -824 -1393 -811
rect -1811 -825 -1623 -824
rect -1581 -825 -1393 -824
rect -1811 -837 -1810 -825
tri -1810 -829 -1806 -825 ne
tri -1398 -829 -1394 -825 nw
rect -1394 -837 -1393 -825
rect -811 -824 -810 -811
tri -810 -824 -806 -820 se
tri -398 -824 -394 -820 sw
rect -394 -824 -393 -811
rect -811 -825 -623 -824
rect -581 -825 -393 -824
rect -811 -837 -810 -825
tri -810 -829 -806 -825 ne
tri -398 -829 -394 -825 nw
rect -394 -837 -393 -825
rect 189 -824 190 -811
tri 190 -824 194 -820 se
tri 602 -824 606 -820 sw
rect 606 -824 607 -811
rect 189 -825 377 -824
rect 419 -825 607 -824
rect 189 -837 190 -825
tri 190 -829 194 -825 ne
tri 602 -829 606 -825 nw
rect 606 -837 607 -825
rect 1189 -824 1190 -811
tri 1190 -824 1194 -820 se
tri 1602 -824 1606 -820 sw
rect 1606 -824 1607 -811
rect 1189 -825 1377 -824
rect 1419 -825 1607 -824
rect 1189 -837 1190 -825
tri 1190 -829 1194 -825 ne
tri 1602 -829 1606 -825 nw
rect 1606 -837 1607 -825
rect 2189 -824 2190 -811
tri 2190 -824 2194 -820 se
tri 2602 -824 2606 -820 sw
rect 2606 -824 2607 -811
rect 2189 -825 2377 -824
rect 2419 -825 2607 -824
rect 2189 -837 2190 -825
tri 2190 -829 2194 -825 ne
tri 2602 -829 2606 -825 nw
rect 2606 -837 2607 -825
rect 3189 -824 3190 -811
tri 3190 -824 3194 -820 se
tri 3602 -824 3606 -820 sw
rect 3606 -824 3607 -811
rect 3189 -825 3377 -824
rect 3419 -825 3607 -824
rect 3189 -837 3190 -825
tri 3190 -829 3194 -825 ne
tri 3602 -829 3606 -825 nw
rect 3606 -837 3607 -825
rect -3638 -864 -3637 -851
tri -3637 -864 -3633 -860 se
tri -3571 -864 -3567 -860 sw
rect -3567 -864 -3566 -851
rect -3638 -865 -3566 -864
rect -3638 -877 -3637 -865
tri -3637 -869 -3633 -865 ne
tri -3571 -869 -3567 -865 nw
rect -3567 -877 -3566 -865
rect -2638 -864 -2637 -851
tri -2637 -864 -2633 -860 se
tri -2571 -864 -2567 -860 sw
rect -2567 -864 -2566 -851
rect -2638 -865 -2566 -864
rect -2638 -877 -2637 -865
tri -2637 -869 -2633 -865 ne
tri -2571 -869 -2567 -865 nw
rect -2567 -877 -2566 -865
rect -1638 -864 -1637 -851
tri -1637 -864 -1633 -860 se
tri -1571 -864 -1567 -860 sw
rect -1567 -864 -1566 -851
rect -1638 -865 -1566 -864
rect -1638 -877 -1637 -865
tri -1637 -869 -1633 -865 ne
tri -1571 -869 -1567 -865 nw
rect -1567 -877 -1566 -865
rect -638 -864 -637 -851
tri -637 -864 -633 -860 se
tri -571 -864 -567 -860 sw
rect -567 -864 -566 -851
rect -638 -865 -566 -864
rect -638 -877 -637 -865
tri -637 -869 -633 -865 ne
tri -571 -869 -567 -865 nw
rect -567 -877 -566 -865
rect 362 -864 363 -851
tri 363 -864 367 -860 se
tri 429 -864 433 -860 sw
rect 433 -864 434 -851
rect 362 -865 434 -864
rect 362 -877 363 -865
tri 363 -869 367 -865 ne
tri 429 -869 433 -865 nw
rect 433 -877 434 -865
rect 1362 -864 1363 -851
tri 1363 -864 1367 -860 se
tri 1429 -864 1433 -860 sw
rect 1433 -864 1434 -851
rect 1362 -865 1434 -864
rect 1362 -877 1363 -865
tri 1363 -869 1367 -865 ne
tri 1429 -869 1433 -865 nw
rect 1433 -877 1434 -865
rect 2362 -864 2363 -851
tri 2363 -864 2367 -860 se
tri 2429 -864 2433 -860 sw
rect 2433 -864 2434 -851
rect 2362 -865 2434 -864
rect 2362 -877 2363 -865
tri 2363 -869 2367 -865 ne
tri 2429 -869 2433 -865 nw
rect 2433 -877 2434 -865
rect 3362 -864 3363 -851
tri 3363 -864 3367 -860 se
tri 3429 -864 3433 -860 sw
rect 3433 -864 3434 -851
rect 3362 -865 3434 -864
rect 3362 -877 3363 -865
tri 3363 -869 3367 -865 ne
tri 3429 -869 3433 -865 nw
rect 3433 -877 3434 -865
rect -974 -1217 -973 -1204
tri -973 -1217 -969 -1213 se
tri -235 -1217 -231 -1213 sw
rect -231 -1217 -230 -1204
rect -974 -1218 -629 -1217
rect -576 -1218 -230 -1217
rect -974 -1230 -973 -1218
tri -973 -1222 -969 -1218 ne
tri -235 -1222 -231 -1218 nw
rect -231 -1230 -230 -1218
rect 26 -1217 27 -1204
tri 27 -1217 31 -1213 se
tri 765 -1217 769 -1213 sw
rect 769 -1217 770 -1204
rect 26 -1218 371 -1217
rect 424 -1218 770 -1217
rect 26 -1230 27 -1218
tri 27 -1222 31 -1218 ne
tri 765 -1222 769 -1218 nw
rect 769 -1230 770 -1218
rect 1026 -1217 1027 -1204
tri 1027 -1217 1031 -1213 se
tri 1765 -1217 1769 -1213 sw
rect 1769 -1217 1770 -1204
rect 1026 -1218 1371 -1217
rect 1424 -1218 1770 -1217
rect 1026 -1230 1027 -1218
tri 1027 -1222 1031 -1218 ne
tri 1765 -1222 1769 -1218 nw
rect 1769 -1230 1770 -1218
rect 2026 -1217 2027 -1204
tri 2027 -1217 2031 -1213 se
tri 2765 -1217 2769 -1213 sw
rect 2769 -1217 2770 -1204
rect 2026 -1218 2371 -1217
rect 2424 -1218 2770 -1217
rect 2026 -1230 2027 -1218
tri 2027 -1222 2031 -1218 ne
tri 2765 -1222 2769 -1218 nw
rect 2769 -1230 2770 -1218
rect 3026 -1217 3027 -1204
tri 3027 -1217 3031 -1213 se
tri 3765 -1217 3769 -1213 sw
rect 3769 -1217 3770 -1204
rect 3026 -1218 3371 -1217
rect 3424 -1218 3770 -1217
rect 3026 -1230 3027 -1218
tri 3027 -1222 3031 -1218 ne
tri 3765 -1222 3769 -1218 nw
rect 3769 -1230 3770 -1218
rect -847 -1380 -846 -1367
tri -846 -1380 -842 -1376 se
tri -362 -1380 -358 -1376 sw
rect -358 -1380 -357 -1367
rect -847 -1381 -655 -1380
rect -548 -1381 -357 -1380
rect -847 -1393 -846 -1381
tri -846 -1385 -842 -1381 ne
tri -362 -1385 -358 -1381 nw
rect -358 -1393 -357 -1381
rect 153 -1380 154 -1367
tri 154 -1380 158 -1376 se
tri 638 -1380 642 -1376 sw
rect 642 -1380 643 -1367
rect 153 -1381 345 -1380
rect 452 -1381 643 -1380
rect 153 -1393 154 -1381
tri 154 -1385 158 -1381 ne
tri 638 -1385 642 -1381 nw
rect 642 -1393 643 -1381
rect 1153 -1380 1154 -1367
tri 1154 -1380 1158 -1376 se
tri 1638 -1380 1642 -1376 sw
rect 1642 -1380 1643 -1367
rect 1153 -1381 1345 -1380
rect 1452 -1381 1643 -1380
rect 1153 -1393 1154 -1381
tri 1154 -1385 1158 -1381 ne
tri 1638 -1385 1642 -1381 nw
rect 1642 -1393 1643 -1381
rect 2153 -1380 2154 -1367
tri 2154 -1380 2158 -1376 se
tri 2638 -1380 2642 -1376 sw
rect 2642 -1380 2643 -1367
rect 2153 -1381 2345 -1380
rect 2452 -1381 2643 -1380
rect 2153 -1393 2154 -1381
tri 2154 -1385 2158 -1381 ne
tri 2638 -1385 2642 -1381 nw
rect 2642 -1393 2643 -1381
rect 3153 -1380 3154 -1367
tri 3154 -1380 3158 -1376 se
tri 3638 -1380 3642 -1376 sw
rect 3642 -1380 3643 -1367
rect 3153 -1381 3345 -1380
rect 3452 -1381 3643 -1380
rect 3153 -1393 3154 -1381
tri 3154 -1385 3158 -1381 ne
tri 3638 -1385 3642 -1381 nw
rect 3642 -1393 3643 -1381
rect -811 -1435 -810 -1422
tri -810 -1435 -806 -1431 se
tri -792 -1435 -788 -1431 sw
rect -788 -1435 -787 -1422
rect -811 -1436 -787 -1435
rect -811 -1448 -810 -1436
tri -810 -1440 -806 -1436 ne
tri -801 -1440 -799 -1437 se
tri -792 -1440 -788 -1436 nw
tri -802 -1443 -801 -1440 se
rect -801 -1443 -799 -1440
tri -799 -1443 -798 -1440 sw
rect -803 -1444 -802 -1443
tri -802 -1444 -801 -1443 nw
rect -799 -1444 -798 -1443
rect -805 -1476 -800 -1444
rect -788 -1448 -787 -1436
rect 189 -1435 190 -1422
tri 190 -1435 194 -1431 se
tri 208 -1435 212 -1431 sw
rect 212 -1435 213 -1422
rect 189 -1436 213 -1435
rect 189 -1448 190 -1436
tri 190 -1440 194 -1436 ne
tri 199 -1440 201 -1437 se
tri 198 -1443 199 -1440 se
rect 199 -1443 201 -1440
tri 201 -1443 202 -1437 sw
tri 208 -1440 212 -1436 nw
rect 197 -1444 198 -1443
tri 198 -1444 199 -1443 nw
rect 201 -1444 202 -1443
rect -393 -1467 -392 -1454
tri -392 -1467 -388 -1463 se
tri -336 -1467 -332 -1463 sw
rect -332 -1467 -331 -1454
rect -393 -1468 -331 -1467
rect -393 -1480 -392 -1468
tri -392 -1472 -388 -1468 ne
tri -336 -1472 -332 -1468 nw
rect -332 -1480 -331 -1468
rect 195 -1476 200 -1444
rect 212 -1448 213 -1436
rect 1189 -1435 1190 -1422
tri 1190 -1435 1194 -1431 se
tri 1208 -1435 1212 -1431 sw
rect 1212 -1435 1213 -1422
rect 1189 -1436 1213 -1435
rect 1189 -1448 1190 -1436
tri 1190 -1440 1194 -1436 ne
tri 1199 -1440 1201 -1437 se
tri 1208 -1440 1212 -1436 nw
tri 1198 -1443 1199 -1440 se
rect 1199 -1443 1201 -1440
tri 1201 -1443 1202 -1440 sw
rect 1197 -1444 1198 -1443
tri 1198 -1444 1199 -1443 nw
rect 1201 -1444 1202 -1443
rect 607 -1467 608 -1454
tri 608 -1467 612 -1463 se
tri 664 -1467 668 -1463 sw
rect 668 -1467 669 -1454
rect 607 -1468 669 -1467
rect 607 -1480 608 -1468
tri 608 -1472 612 -1468 ne
tri 664 -1472 668 -1468 nw
rect 668 -1480 669 -1468
rect 1195 -1476 1200 -1444
rect 1212 -1448 1213 -1436
rect 2189 -1435 2190 -1422
tri 2190 -1435 2194 -1431 se
tri 2208 -1435 2212 -1431 sw
rect 2212 -1435 2213 -1422
rect 2189 -1436 2213 -1435
rect 2189 -1448 2190 -1436
tri 2190 -1440 2194 -1436 ne
tri 2199 -1440 2201 -1437 se
tri 2208 -1440 2212 -1436 nw
tri 2198 -1443 2199 -1440 se
rect 2199 -1443 2201 -1440
tri 2201 -1443 2202 -1440 sw
rect 2197 -1444 2198 -1443
tri 2198 -1444 2199 -1443 nw
rect 2201 -1444 2202 -1443
rect 1607 -1467 1608 -1454
tri 1608 -1467 1612 -1463 se
tri 1664 -1467 1668 -1463 sw
rect 1668 -1467 1669 -1454
rect 1607 -1468 1669 -1467
rect 1607 -1480 1608 -1468
tri 1608 -1472 1612 -1468 ne
tri 1664 -1472 1668 -1468 nw
rect 1668 -1480 1669 -1468
rect 2195 -1476 2200 -1444
rect 2212 -1448 2213 -1436
rect 3189 -1435 3190 -1422
tri 3190 -1435 3194 -1431 se
tri 3208 -1435 3212 -1431 sw
rect 3212 -1435 3213 -1422
rect 3189 -1436 3213 -1435
rect 3189 -1448 3190 -1436
tri 3190 -1440 3194 -1436 ne
tri 3199 -1440 3201 -1437 se
tri 3208 -1440 3212 -1436 nw
tri 3198 -1443 3199 -1440 se
rect 3199 -1443 3201 -1440
tri 3201 -1443 3202 -1440 sw
rect 3197 -1444 3198 -1443
tri 3198 -1444 3199 -1443 nw
rect 3201 -1444 3202 -1443
rect 2607 -1467 2608 -1454
tri 2608 -1467 2612 -1463 se
tri 2664 -1467 2668 -1463 sw
rect 2668 -1467 2669 -1454
rect 2607 -1468 2669 -1467
rect 2607 -1480 2608 -1468
tri 2608 -1472 2612 -1468 ne
tri 2664 -1472 2668 -1468 nw
rect 2668 -1480 2669 -1468
rect 3195 -1476 3200 -1444
rect 3212 -1448 3213 -1436
rect 3607 -1467 3608 -1454
tri 3608 -1467 3612 -1463 se
tri 3664 -1467 3668 -1463 sw
rect 3668 -1467 3669 -1454
rect 3607 -1468 3669 -1467
rect 3607 -1480 3608 -1468
tri 3608 -1472 3612 -1468 ne
tri 3664 -1472 3668 -1468 nw
rect 3668 -1480 3669 -1468
rect -670 -1521 -669 -1508
tri -669 -1521 -665 -1517 se
tri -539 -1521 -535 -1517 sw
rect -535 -1521 -534 -1508
rect -670 -1522 -623 -1521
rect -581 -1522 -534 -1521
rect -670 -1534 -669 -1522
tri -669 -1526 -665 -1522 ne
tri -539 -1526 -535 -1522 nw
rect -535 -1534 -534 -1522
rect 330 -1521 331 -1508
tri 331 -1521 335 -1517 se
tri 461 -1521 465 -1517 sw
rect 465 -1521 466 -1508
rect 330 -1522 377 -1521
rect 419 -1522 466 -1521
rect 330 -1534 331 -1522
tri 331 -1526 335 -1522 ne
tri 461 -1526 465 -1522 nw
rect 465 -1534 466 -1522
rect 1330 -1521 1331 -1508
tri 1331 -1521 1335 -1517 se
tri 1461 -1521 1465 -1517 sw
rect 1465 -1521 1466 -1508
rect 1330 -1522 1377 -1521
rect 1419 -1522 1466 -1521
rect 1330 -1534 1331 -1522
tri 1331 -1526 1335 -1522 ne
tri 1461 -1526 1465 -1522 nw
rect 1465 -1534 1466 -1522
rect 2330 -1521 2331 -1508
tri 2331 -1521 2335 -1517 se
tri 2461 -1521 2465 -1517 sw
rect 2465 -1521 2466 -1508
rect 2330 -1522 2377 -1521
rect 2419 -1522 2466 -1521
rect 2330 -1534 2331 -1522
tri 2331 -1526 2335 -1522 ne
tri 2461 -1526 2465 -1522 nw
rect 2465 -1534 2466 -1522
rect 3330 -1521 3331 -1508
tri 3331 -1521 3335 -1517 se
tri 3461 -1521 3465 -1517 sw
rect 3465 -1521 3466 -1508
rect 3330 -1522 3377 -1521
rect 3419 -1522 3466 -1521
rect 3330 -1534 3331 -1522
tri 3331 -1526 3335 -1522 ne
tri 3461 -1526 3465 -1522 nw
rect 3465 -1534 3466 -1522
rect -811 -1558 -810 -1545
tri -810 -1558 -806 -1554 se
tri -744 -1558 -740 -1554 sw
rect -740 -1558 -739 -1545
rect -811 -1559 -739 -1558
rect -811 -1571 -810 -1559
tri -810 -1563 -806 -1559 ne
tri -744 -1563 -740 -1559 nw
rect -740 -1571 -739 -1559
rect 189 -1558 190 -1545
tri 190 -1558 194 -1554 se
tri 256 -1558 260 -1554 sw
rect 260 -1558 261 -1545
rect 189 -1559 261 -1558
rect 189 -1571 190 -1559
tri 190 -1563 194 -1559 ne
tri 256 -1563 260 -1559 nw
rect 260 -1571 261 -1559
rect 1189 -1558 1190 -1545
tri 1190 -1558 1194 -1554 se
tri 1256 -1558 1260 -1554 sw
rect 1260 -1558 1261 -1545
rect 1189 -1559 1261 -1558
rect 1189 -1571 1190 -1559
tri 1190 -1563 1194 -1559 ne
tri 1256 -1563 1260 -1559 nw
rect 1260 -1571 1261 -1559
rect 2189 -1558 2190 -1545
tri 2190 -1558 2194 -1554 se
tri 2256 -1558 2260 -1554 sw
rect 2260 -1558 2261 -1545
rect 2189 -1559 2261 -1558
rect 2189 -1571 2190 -1559
tri 2190 -1563 2194 -1559 ne
tri 2256 -1563 2260 -1559 nw
rect 2260 -1571 2261 -1559
rect 3189 -1558 3190 -1545
tri 3190 -1558 3194 -1554 se
tri 3256 -1558 3260 -1554 sw
rect 3260 -1558 3261 -1545
rect 3189 -1559 3261 -1558
rect 3189 -1571 3190 -1559
tri 3190 -1563 3194 -1559 ne
tri 3256 -1563 3260 -1559 nw
rect 3260 -1571 3261 -1559
tri -610 -1596 -608 -1594 se
tri -608 -1596 -607 -1594 sw
tri -597 -1596 -596 -1594 se
tri -596 -1596 -594 -1594 sw
tri -610 -1597 -608 -1596 ne
rect -608 -1597 -607 -1596
tri -607 -1597 -605 -1596 sw
tri -599 -1597 -597 -1596 se
tri -608 -1600 -605 -1597 ne
tri -605 -1599 -604 -1597 sw
tri -600 -1599 -599 -1597 se
rect -599 -1599 -597 -1597
tri -597 -1599 -594 -1596 nw
tri 390 -1596 392 -1594 se
tri 392 -1596 393 -1594 sw
tri 403 -1596 404 -1594 se
tri 404 -1596 406 -1594 sw
tri 390 -1597 392 -1596 ne
rect 392 -1597 393 -1596
tri 393 -1597 395 -1596 sw
tri 401 -1597 403 -1596 se
rect -605 -1600 -604 -1599
tri -604 -1600 -602 -1599 sw
tri -602 -1600 -600 -1599 se
tri -605 -1602 -604 -1600 ne
tri -607 -1605 -604 -1602 se
rect -604 -1604 -600 -1600
tri -600 -1602 -597 -1599 nw
tri 392 -1600 395 -1597 ne
tri 395 -1599 396 -1597 sw
tri 400 -1599 401 -1597 se
rect 401 -1599 403 -1597
tri 403 -1599 406 -1596 nw
tri 1390 -1596 1392 -1594 se
tri 1392 -1596 1393 -1594 sw
tri 1403 -1596 1404 -1594 se
tri 1404 -1596 1406 -1594 sw
tri 1390 -1597 1392 -1596 ne
rect 1392 -1597 1393 -1596
tri 1393 -1597 1395 -1596 sw
tri 1401 -1597 1403 -1596 se
rect 395 -1600 396 -1599
tri 396 -1600 398 -1599 sw
tri 398 -1600 400 -1599 se
tri 395 -1602 396 -1600 ne
rect -604 -1605 -603 -1604
tri -603 -1605 -602 -1604 nw
tri -602 -1605 -601 -1604 ne
rect -601 -1605 -600 -1604
tri -600 -1605 -597 -1602 sw
tri 393 -1605 396 -1602 se
rect 396 -1604 400 -1600
tri 400 -1602 403 -1599 nw
tri 1392 -1600 1395 -1597 ne
tri 1395 -1599 1396 -1597 sw
tri 1400 -1599 1401 -1597 se
rect 1401 -1599 1403 -1597
tri 1403 -1599 1406 -1596 nw
tri 2390 -1596 2392 -1594 se
tri 2392 -1596 2393 -1594 sw
tri 2403 -1596 2404 -1594 se
tri 2404 -1596 2406 -1594 sw
tri 2390 -1597 2392 -1596 ne
rect 2392 -1597 2393 -1596
tri 2393 -1597 2395 -1596 sw
tri 2401 -1597 2403 -1596 se
rect 1395 -1600 1396 -1599
tri 1396 -1600 1398 -1599 sw
tri 1398 -1600 1400 -1599 se
tri 1395 -1602 1396 -1600 ne
rect 396 -1605 397 -1604
tri 397 -1605 398 -1604 nw
tri 398 -1605 399 -1604 ne
rect 399 -1605 400 -1604
tri 400 -1605 403 -1602 sw
tri 1393 -1605 1396 -1602 se
rect 1396 -1604 1400 -1600
tri 1400 -1602 1403 -1599 nw
tri 2392 -1600 2395 -1597 ne
tri 2395 -1599 2396 -1597 sw
tri 2400 -1599 2401 -1597 se
rect 2401 -1599 2403 -1597
tri 2403 -1599 2406 -1596 nw
tri 3390 -1596 3392 -1594 se
tri 3392 -1596 3393 -1594 sw
tri 3403 -1596 3404 -1594 se
tri 3404 -1596 3406 -1594 sw
tri 3390 -1597 3392 -1596 ne
rect 3392 -1597 3393 -1596
tri 3393 -1597 3395 -1596 sw
tri 3401 -1597 3403 -1596 se
rect 2395 -1600 2396 -1599
tri 2396 -1600 2398 -1599 sw
tri 2398 -1600 2400 -1599 se
tri 2395 -1602 2396 -1600 ne
rect 1396 -1605 1397 -1604
tri 1397 -1605 1398 -1604 nw
tri 1398 -1605 1399 -1604 ne
rect 1399 -1605 1400 -1604
tri 1400 -1605 1403 -1602 sw
tri 2393 -1605 2396 -1602 se
rect 2396 -1604 2400 -1600
tri 2400 -1602 2403 -1599 nw
tri 3392 -1600 3395 -1597 ne
tri 3395 -1599 3396 -1597 sw
tri 3400 -1599 3401 -1597 se
rect 3401 -1599 3403 -1597
tri 3403 -1599 3406 -1596 nw
rect 3395 -1600 3396 -1599
tri 3396 -1600 3398 -1599 sw
tri 3398 -1600 3400 -1599 se
tri 3395 -1602 3396 -1600 ne
rect 2396 -1605 2397 -1604
tri 2397 -1605 2398 -1604 nw
tri 2398 -1605 2399 -1604 ne
rect 2399 -1605 2400 -1604
tri 2400 -1605 2403 -1602 sw
tri 3393 -1605 3396 -1602 se
rect 3396 -1604 3400 -1600
tri 3400 -1602 3403 -1599 nw
rect 3396 -1605 3397 -1604
tri 3397 -1605 3398 -1604 nw
tri 3398 -1605 3399 -1604 ne
rect 3399 -1605 3400 -1604
tri 3400 -1605 3403 -1602 sw
tri -610 -1608 -607 -1605 se
tri -607 -1608 -604 -1605 nw
tri -600 -1608 -597 -1605 ne
tri -597 -1608 -594 -1605 sw
tri -610 -1610 -608 -1608 ne
tri -608 -1610 -607 -1608 nw
tri -597 -1610 -596 -1608 ne
tri -596 -1610 -594 -1608 nw
tri 390 -1608 393 -1605 se
tri 393 -1608 396 -1605 nw
tri 400 -1608 403 -1605 ne
tri 403 -1608 406 -1605 sw
tri 390 -1610 392 -1608 ne
tri 392 -1610 393 -1608 nw
tri 403 -1610 404 -1608 ne
tri 404 -1610 406 -1608 nw
tri 1390 -1608 1393 -1605 se
tri 1393 -1608 1396 -1605 nw
tri 1400 -1608 1403 -1605 ne
tri 1403 -1608 1406 -1605 sw
tri 1390 -1610 1392 -1608 ne
tri 1392 -1610 1393 -1608 nw
tri 1403 -1610 1404 -1608 ne
tri 1404 -1610 1406 -1608 nw
tri 2390 -1608 2393 -1605 se
tri 2393 -1608 2396 -1605 nw
tri 2400 -1608 2403 -1605 ne
tri 2403 -1608 2406 -1605 sw
tri 2390 -1610 2392 -1608 ne
tri 2392 -1610 2393 -1608 nw
tri 2403 -1610 2404 -1608 ne
tri 2404 -1610 2406 -1608 nw
tri 3390 -1608 3393 -1605 se
tri 3393 -1608 3396 -1605 nw
tri 3400 -1608 3403 -1605 ne
tri 3403 -1608 3406 -1605 sw
tri 3390 -1610 3392 -1608 ne
tri 3392 -1610 3393 -1608 nw
tri 3403 -1610 3404 -1608 ne
tri 3404 -1610 3406 -1608 nw
rect -534 -1670 -533 -1657
tri -533 -1670 -529 -1666 se
tri -470 -1670 -466 -1666 sw
rect -466 -1670 -465 -1657
rect -534 -1671 -465 -1670
rect -534 -1683 -533 -1671
tri -533 -1675 -529 -1671 ne
tri -470 -1675 -466 -1671 nw
rect -466 -1683 -465 -1671
rect -331 -1670 -330 -1657
tri -330 -1670 -326 -1666 se
tri -235 -1670 -231 -1666 sw
rect -231 -1670 -230 -1657
rect -331 -1671 -230 -1670
rect -331 -1683 -330 -1671
tri -330 -1675 -326 -1671 ne
tri -235 -1675 -231 -1671 nw
rect -231 -1683 -230 -1671
rect 466 -1670 467 -1657
tri 467 -1670 471 -1666 se
tri 530 -1670 534 -1666 sw
rect 534 -1670 535 -1657
rect 466 -1671 535 -1670
rect 466 -1683 467 -1671
tri 467 -1675 471 -1671 ne
tri 530 -1675 534 -1671 nw
rect 534 -1683 535 -1671
rect 669 -1670 670 -1657
tri 670 -1670 674 -1666 se
tri 765 -1670 769 -1666 sw
rect 769 -1670 770 -1657
rect 669 -1671 770 -1670
rect 669 -1683 670 -1671
tri 670 -1675 674 -1671 ne
tri 765 -1675 769 -1671 nw
rect 769 -1683 770 -1671
rect 1466 -1670 1467 -1657
tri 1467 -1670 1471 -1666 se
tri 1530 -1670 1534 -1666 sw
rect 1534 -1670 1535 -1657
rect 1466 -1671 1535 -1670
rect 1466 -1683 1467 -1671
tri 1467 -1675 1471 -1671 ne
tri 1530 -1675 1534 -1671 nw
rect 1534 -1683 1535 -1671
rect 1669 -1670 1670 -1657
tri 1670 -1670 1674 -1666 se
tri 1765 -1670 1769 -1666 sw
rect 1769 -1670 1770 -1657
rect 1669 -1671 1770 -1670
rect 1669 -1683 1670 -1671
tri 1670 -1675 1674 -1671 ne
tri 1765 -1675 1769 -1671 nw
rect 1769 -1683 1770 -1671
rect 2466 -1670 2467 -1657
tri 2467 -1670 2471 -1666 se
tri 2530 -1670 2534 -1666 sw
rect 2534 -1670 2535 -1657
rect 2466 -1671 2535 -1670
rect 2466 -1683 2467 -1671
tri 2467 -1675 2471 -1671 ne
tri 2530 -1675 2534 -1671 nw
rect 2534 -1683 2535 -1671
rect 2669 -1670 2670 -1657
tri 2670 -1670 2674 -1666 se
tri 2765 -1670 2769 -1666 sw
rect 2769 -1670 2770 -1657
rect 2669 -1671 2770 -1670
rect 2669 -1683 2670 -1671
tri 2670 -1675 2674 -1671 ne
tri 2765 -1675 2769 -1671 nw
rect 2769 -1683 2770 -1671
rect 3466 -1670 3467 -1657
tri 3467 -1670 3471 -1666 se
tri 3530 -1670 3534 -1666 sw
rect 3534 -1670 3535 -1657
rect 3466 -1671 3535 -1670
rect 3466 -1683 3467 -1671
tri 3467 -1675 3471 -1671 ne
tri 3530 -1675 3534 -1671 nw
rect 3534 -1683 3535 -1671
rect 3669 -1670 3670 -1657
tri 3670 -1670 3674 -1666 se
tri 3765 -1670 3769 -1666 sw
rect 3769 -1670 3770 -1657
rect 3669 -1671 3770 -1670
rect 3669 -1683 3670 -1671
tri 3670 -1675 3674 -1671 ne
tri 3765 -1675 3769 -1671 nw
rect 3769 -1683 3770 -1671
rect -811 -1824 -810 -1811
tri -810 -1824 -806 -1820 se
tri -398 -1824 -394 -1820 sw
rect -394 -1824 -393 -1811
rect -811 -1825 -623 -1824
rect -581 -1825 -393 -1824
rect -811 -1837 -810 -1825
tri -810 -1829 -806 -1825 ne
tri -398 -1829 -394 -1825 nw
rect -394 -1837 -393 -1825
rect 189 -1824 190 -1811
tri 190 -1824 194 -1820 se
tri 602 -1824 606 -1820 sw
rect 606 -1824 607 -1811
rect 189 -1825 377 -1824
rect 419 -1825 607 -1824
rect 189 -1837 190 -1825
tri 190 -1829 194 -1825 ne
tri 602 -1829 606 -1825 nw
rect 606 -1837 607 -1825
rect 1189 -1824 1190 -1811
tri 1190 -1824 1194 -1820 se
tri 1602 -1824 1606 -1820 sw
rect 1606 -1824 1607 -1811
rect 1189 -1825 1377 -1824
rect 1419 -1825 1607 -1824
rect 1189 -1837 1190 -1825
tri 1190 -1829 1194 -1825 ne
tri 1602 -1829 1606 -1825 nw
rect 1606 -1837 1607 -1825
rect 2189 -1824 2190 -1811
tri 2190 -1824 2194 -1820 se
tri 2602 -1824 2606 -1820 sw
rect 2606 -1824 2607 -1811
rect 2189 -1825 2377 -1824
rect 2419 -1825 2607 -1824
rect 2189 -1837 2190 -1825
tri 2190 -1829 2194 -1825 ne
tri 2602 -1829 2606 -1825 nw
rect 2606 -1837 2607 -1825
rect 3189 -1824 3190 -1811
tri 3190 -1824 3194 -1820 se
tri 3602 -1824 3606 -1820 sw
rect 3606 -1824 3607 -1811
rect 3189 -1825 3377 -1824
rect 3419 -1825 3607 -1824
rect 3189 -1837 3190 -1825
tri 3190 -1829 3194 -1825 ne
tri 3602 -1829 3606 -1825 nw
rect 3606 -1837 3607 -1825
rect -638 -1864 -637 -1851
tri -637 -1864 -633 -1860 se
tri -571 -1864 -567 -1860 sw
rect -567 -1864 -566 -1851
rect -638 -1865 -566 -1864
rect -638 -1877 -637 -1865
tri -637 -1869 -633 -1865 ne
tri -571 -1869 -567 -1865 nw
rect -567 -1877 -566 -1865
rect 362 -1864 363 -1851
tri 363 -1864 367 -1860 se
tri 429 -1864 433 -1860 sw
rect 433 -1864 434 -1851
rect 362 -1865 434 -1864
rect 362 -1877 363 -1865
tri 363 -1869 367 -1865 ne
tri 429 -1869 433 -1865 nw
rect 433 -1877 434 -1865
rect 1362 -1864 1363 -1851
tri 1363 -1864 1367 -1860 se
tri 1429 -1864 1433 -1860 sw
rect 1433 -1864 1434 -1851
rect 1362 -1865 1434 -1864
rect 1362 -1877 1363 -1865
tri 1363 -1869 1367 -1865 ne
tri 1429 -1869 1433 -1865 nw
rect 1433 -1877 1434 -1865
rect 2362 -1864 2363 -1851
tri 2363 -1864 2367 -1860 se
tri 2429 -1864 2433 -1860 sw
rect 2433 -1864 2434 -1851
rect 2362 -1865 2434 -1864
rect 2362 -1877 2363 -1865
tri 2363 -1869 2367 -1865 ne
tri 2429 -1869 2433 -1865 nw
rect 2433 -1877 2434 -1865
rect 3362 -1864 3363 -1851
tri 3363 -1864 3367 -1860 se
tri 3429 -1864 3433 -1860 sw
rect 3433 -1864 3434 -1851
rect 3362 -1865 3434 -1864
rect 3362 -1877 3363 -1865
tri 3363 -1869 3367 -1865 ne
tri 3429 -1869 3433 -1865 nw
rect 3433 -1877 3434 -1865
rect -974 -2217 -973 -2204
tri -973 -2217 -969 -2213 se
tri -235 -2217 -231 -2213 sw
rect -231 -2217 -230 -2204
rect -974 -2218 -629 -2217
rect -576 -2218 -230 -2217
rect -974 -2230 -973 -2218
tri -973 -2222 -969 -2218 ne
tri -235 -2222 -231 -2218 nw
rect -231 -2230 -230 -2218
rect 26 -2217 27 -2204
tri 27 -2217 31 -2213 se
tri 765 -2217 769 -2213 sw
rect 769 -2217 770 -2204
rect 26 -2218 371 -2217
rect 424 -2218 770 -2217
rect 26 -2230 27 -2218
tri 27 -2222 31 -2218 ne
tri 765 -2222 769 -2218 nw
rect 769 -2230 770 -2218
rect 1026 -2217 1027 -2204
tri 1027 -2217 1031 -2213 se
tri 1765 -2217 1769 -2213 sw
rect 1769 -2217 1770 -2204
rect 1026 -2218 1371 -2217
rect 1424 -2218 1770 -2217
rect 1026 -2230 1027 -2218
tri 1027 -2222 1031 -2218 ne
tri 1765 -2222 1769 -2218 nw
rect 1769 -2230 1770 -2218
rect 2026 -2217 2027 -2204
tri 2027 -2217 2031 -2213 se
tri 2765 -2217 2769 -2213 sw
rect 2769 -2217 2770 -2204
rect 2026 -2218 2371 -2217
rect 2424 -2218 2770 -2217
rect 2026 -2230 2027 -2218
tri 2027 -2222 2031 -2218 ne
tri 2765 -2222 2769 -2218 nw
rect 2769 -2230 2770 -2218
rect 3026 -2217 3027 -2204
tri 3027 -2217 3031 -2213 se
tri 3765 -2217 3769 -2213 sw
rect 3769 -2217 3770 -2204
rect 3026 -2218 3371 -2217
rect 3424 -2218 3770 -2217
rect 3026 -2230 3027 -2218
tri 3027 -2222 3031 -2218 ne
tri 3765 -2222 3769 -2218 nw
rect 3769 -2230 3770 -2218
rect -847 -2380 -846 -2367
tri -846 -2380 -842 -2376 se
tri -362 -2380 -358 -2376 sw
rect -358 -2380 -357 -2367
rect -847 -2381 -655 -2380
rect -548 -2381 -357 -2380
rect -847 -2393 -846 -2381
tri -846 -2385 -842 -2381 ne
tri -362 -2385 -358 -2381 nw
rect -358 -2393 -357 -2381
rect 153 -2380 154 -2367
tri 154 -2380 158 -2376 se
tri 638 -2380 642 -2376 sw
rect 642 -2380 643 -2367
rect 153 -2381 345 -2380
rect 452 -2381 643 -2380
rect 153 -2393 154 -2381
tri 154 -2385 158 -2381 ne
tri 638 -2385 642 -2381 nw
rect 642 -2393 643 -2381
rect 1153 -2380 1154 -2367
tri 1154 -2380 1158 -2376 se
tri 1638 -2380 1642 -2376 sw
rect 1642 -2380 1643 -2367
rect 1153 -2381 1345 -2380
rect 1452 -2381 1643 -2380
rect 1153 -2393 1154 -2381
tri 1154 -2385 1158 -2381 ne
tri 1638 -2385 1642 -2381 nw
rect 1642 -2393 1643 -2381
rect 2153 -2380 2154 -2367
tri 2154 -2380 2158 -2376 se
tri 2638 -2380 2642 -2376 sw
rect 2642 -2380 2643 -2367
rect 2153 -2381 2345 -2380
rect 2452 -2381 2643 -2380
rect 2153 -2393 2154 -2381
tri 2154 -2385 2158 -2381 ne
tri 2638 -2385 2642 -2381 nw
rect 2642 -2393 2643 -2381
rect 3153 -2380 3154 -2367
tri 3154 -2380 3158 -2376 se
tri 3638 -2380 3642 -2376 sw
rect 3642 -2380 3643 -2367
rect 3153 -2381 3345 -2380
rect 3452 -2381 3643 -2380
rect 3153 -2393 3154 -2381
tri 3154 -2385 3158 -2381 ne
tri 3638 -2385 3642 -2381 nw
rect 3642 -2393 3643 -2381
rect -811 -2435 -810 -2422
tri -810 -2435 -806 -2431 se
tri -792 -2435 -788 -2431 sw
rect -788 -2435 -787 -2422
rect -811 -2436 -787 -2435
rect -811 -2448 -810 -2436
tri -810 -2440 -806 -2436 ne
tri -801 -2440 -799 -2437 se
tri -792 -2440 -788 -2436 nw
tri -802 -2443 -801 -2440 se
rect -801 -2443 -799 -2440
tri -799 -2443 -798 -2440 sw
rect -803 -2444 -802 -2443
tri -802 -2444 -801 -2443 nw
rect -799 -2444 -798 -2443
rect -805 -2476 -800 -2444
rect -788 -2448 -787 -2436
rect 189 -2435 190 -2422
tri 190 -2435 194 -2431 se
tri 208 -2435 212 -2431 sw
rect 212 -2435 213 -2422
rect 189 -2436 213 -2435
rect 189 -2448 190 -2436
tri 190 -2440 194 -2436 ne
tri 199 -2440 201 -2437 se
tri 208 -2440 212 -2436 nw
tri 198 -2443 199 -2440 se
rect 199 -2443 201 -2440
tri 201 -2443 202 -2440 sw
rect 197 -2444 198 -2443
tri 198 -2444 199 -2443 nw
rect 201 -2444 202 -2443
rect -393 -2467 -392 -2454
tri -392 -2467 -388 -2463 se
tri -336 -2467 -332 -2463 sw
rect -332 -2467 -331 -2454
rect -393 -2468 -331 -2467
rect -393 -2480 -392 -2468
tri -392 -2472 -388 -2468 ne
tri -336 -2472 -332 -2468 nw
rect -332 -2480 -331 -2468
rect 195 -2476 200 -2444
rect 212 -2448 213 -2436
rect 1189 -2435 1190 -2422
tri 1190 -2435 1194 -2431 se
tri 1208 -2435 1212 -2431 sw
rect 1212 -2435 1213 -2422
rect 1189 -2436 1213 -2435
rect 1189 -2448 1190 -2436
tri 1190 -2440 1194 -2436 ne
tri 1199 -2440 1201 -2437 se
tri 1208 -2440 1212 -2436 nw
tri 1198 -2443 1199 -2440 se
rect 1199 -2443 1201 -2440
tri 1201 -2443 1202 -2440 sw
rect 1197 -2444 1198 -2443
tri 1198 -2444 1199 -2443 nw
rect 1201 -2444 1202 -2443
rect 607 -2467 608 -2454
tri 608 -2467 612 -2463 se
tri 664 -2467 668 -2463 sw
rect 668 -2467 669 -2454
rect 607 -2468 669 -2467
rect 607 -2480 608 -2468
tri 608 -2472 612 -2468 ne
tri 664 -2472 668 -2468 nw
rect 668 -2480 669 -2468
rect 1195 -2476 1200 -2444
rect 1212 -2448 1213 -2436
rect 2189 -2435 2190 -2422
tri 2190 -2435 2194 -2431 se
tri 2208 -2435 2212 -2431 sw
rect 2212 -2435 2213 -2422
rect 2189 -2436 2213 -2435
rect 2189 -2448 2190 -2436
tri 2190 -2440 2194 -2436 ne
tri 2199 -2440 2201 -2437 se
tri 2208 -2440 2212 -2436 nw
tri 2198 -2443 2199 -2440 se
rect 2199 -2443 2201 -2440
tri 2201 -2443 2202 -2440 sw
rect 2197 -2444 2198 -2443
tri 2198 -2444 2199 -2443 nw
rect 2201 -2444 2202 -2443
rect 1607 -2467 1608 -2454
tri 1608 -2467 1612 -2463 se
tri 1664 -2467 1668 -2463 sw
rect 1668 -2467 1669 -2454
rect 1607 -2468 1669 -2467
rect 1607 -2480 1608 -2468
tri 1608 -2472 1612 -2468 ne
tri 1664 -2472 1668 -2468 nw
rect 1668 -2480 1669 -2468
rect 2195 -2476 2200 -2444
rect 2212 -2448 2213 -2436
rect 3189 -2435 3190 -2422
tri 3190 -2435 3194 -2431 se
tri 3208 -2435 3212 -2431 sw
rect 3212 -2435 3213 -2422
rect 3189 -2436 3213 -2435
rect 3189 -2448 3190 -2436
tri 3190 -2440 3194 -2436 ne
tri 3199 -2440 3201 -2437 se
tri 3208 -2440 3212 -2436 nw
tri 3198 -2443 3199 -2440 se
rect 3199 -2443 3201 -2440
tri 3201 -2443 3202 -2440 sw
rect 3197 -2444 3198 -2443
tri 3198 -2444 3199 -2443 nw
rect 3201 -2444 3202 -2443
rect 2607 -2467 2608 -2454
tri 2608 -2467 2612 -2463 se
tri 2664 -2467 2668 -2463 sw
rect 2668 -2467 2669 -2454
rect 2607 -2468 2669 -2467
rect 2607 -2480 2608 -2468
tri 2608 -2472 2612 -2468 ne
tri 2664 -2472 2668 -2468 nw
rect 2668 -2480 2669 -2468
rect 3195 -2476 3200 -2444
rect 3212 -2448 3213 -2436
rect 3607 -2467 3608 -2454
tri 3608 -2467 3612 -2463 se
tri 3664 -2467 3668 -2463 sw
rect 3668 -2467 3669 -2454
rect 3607 -2468 3669 -2467
rect 3607 -2480 3608 -2468
tri 3608 -2472 3612 -2468 ne
tri 3664 -2472 3668 -2468 nw
rect 3668 -2480 3669 -2468
rect -670 -2521 -669 -2508
tri -669 -2521 -665 -2517 se
tri -539 -2521 -535 -2517 sw
rect -535 -2521 -534 -2508
rect -670 -2522 -623 -2521
rect -581 -2522 -534 -2521
rect -670 -2534 -669 -2522
tri -669 -2526 -665 -2522 ne
tri -539 -2526 -535 -2522 nw
rect -535 -2534 -534 -2522
rect 330 -2521 331 -2508
tri 331 -2521 335 -2517 se
tri 461 -2521 465 -2517 sw
rect 465 -2521 466 -2508
rect 330 -2522 377 -2521
rect 419 -2522 466 -2521
rect 330 -2534 331 -2522
tri 331 -2526 335 -2522 ne
tri 461 -2526 465 -2522 nw
rect 465 -2534 466 -2522
rect 1330 -2521 1331 -2508
tri 1331 -2521 1335 -2517 se
tri 1461 -2521 1465 -2517 sw
rect 1465 -2521 1466 -2508
rect 1330 -2522 1377 -2521
rect 1419 -2522 1466 -2521
rect 1330 -2534 1331 -2522
tri 1331 -2526 1335 -2522 ne
tri 1461 -2526 1465 -2522 nw
rect 1465 -2534 1466 -2522
rect 2330 -2521 2331 -2508
tri 2331 -2521 2335 -2517 se
tri 2461 -2521 2465 -2517 sw
rect 2465 -2521 2466 -2508
rect 2330 -2522 2377 -2521
rect 2419 -2522 2466 -2521
rect 2330 -2534 2331 -2522
tri 2331 -2526 2335 -2522 ne
tri 2461 -2526 2465 -2522 nw
rect 2465 -2534 2466 -2522
rect 3330 -2521 3331 -2508
tri 3331 -2521 3335 -2517 se
tri 3461 -2521 3465 -2517 sw
rect 3465 -2521 3466 -2508
rect 3330 -2522 3377 -2521
rect 3419 -2522 3466 -2521
rect 3330 -2534 3331 -2522
tri 3331 -2526 3335 -2522 ne
tri 3461 -2526 3465 -2522 nw
rect 3465 -2534 3466 -2522
rect -811 -2558 -810 -2545
tri -810 -2558 -806 -2554 se
tri -744 -2558 -740 -2554 sw
rect -740 -2558 -739 -2545
rect -811 -2559 -739 -2558
rect -811 -2571 -810 -2559
tri -810 -2563 -806 -2559 ne
tri -744 -2563 -740 -2559 nw
rect -740 -2571 -739 -2559
rect 189 -2558 190 -2545
tri 190 -2558 194 -2554 se
tri 256 -2558 260 -2554 sw
rect 260 -2558 261 -2545
rect 189 -2559 261 -2558
rect 189 -2571 190 -2559
tri 190 -2563 194 -2559 ne
tri 256 -2563 260 -2559 nw
rect 260 -2571 261 -2559
rect 1189 -2558 1190 -2545
tri 1190 -2558 1194 -2554 se
tri 1256 -2558 1260 -2554 sw
rect 1260 -2558 1261 -2545
rect 1189 -2559 1261 -2558
rect 1189 -2571 1190 -2559
tri 1190 -2563 1194 -2559 ne
tri 1256 -2563 1260 -2559 nw
rect 1260 -2571 1261 -2559
rect 2189 -2558 2190 -2545
tri 2190 -2558 2194 -2554 se
tri 2256 -2558 2260 -2554 sw
rect 2260 -2558 2261 -2545
rect 2189 -2559 2261 -2558
rect 2189 -2571 2190 -2559
tri 2190 -2563 2194 -2559 ne
tri 2256 -2563 2260 -2559 nw
rect 2260 -2571 2261 -2559
rect 3189 -2558 3190 -2545
tri 3190 -2558 3194 -2554 se
tri 3256 -2558 3260 -2554 sw
rect 3260 -2558 3261 -2545
rect 3189 -2559 3261 -2558
rect 3189 -2571 3190 -2559
tri 3190 -2563 3194 -2559 ne
tri 3256 -2563 3260 -2559 nw
rect 3260 -2571 3261 -2559
tri -610 -2596 -608 -2594 se
tri -608 -2596 -607 -2594 sw
tri -597 -2596 -596 -2594 se
tri -596 -2596 -594 -2594 sw
tri -610 -2597 -608 -2596 ne
rect -608 -2597 -607 -2596
tri -607 -2597 -605 -2596 sw
tri -599 -2597 -597 -2596 se
tri -608 -2600 -605 -2597 ne
tri -605 -2599 -604 -2597 sw
tri -600 -2599 -599 -2597 se
rect -599 -2599 -597 -2597
tri -597 -2599 -594 -2596 nw
tri 390 -2596 392 -2594 se
tri 392 -2596 393 -2594 sw
tri 403 -2596 404 -2594 se
tri 404 -2596 406 -2594 sw
tri 390 -2597 392 -2596 ne
rect 392 -2597 393 -2596
tri 393 -2597 395 -2596 sw
tri 401 -2597 403 -2596 se
rect -605 -2600 -604 -2599
tri -604 -2600 -602 -2599 sw
tri -602 -2600 -600 -2599 se
tri -605 -2602 -604 -2600 ne
tri -607 -2605 -604 -2602 se
rect -604 -2604 -600 -2600
tri -600 -2602 -597 -2599 nw
tri 392 -2600 395 -2597 ne
tri 395 -2599 396 -2597 sw
tri 400 -2599 401 -2597 se
rect 401 -2599 403 -2597
tri 403 -2599 406 -2596 nw
tri 1390 -2596 1392 -2594 se
tri 1392 -2596 1393 -2594 sw
tri 1403 -2596 1404 -2594 se
tri 1404 -2596 1406 -2594 sw
tri 1390 -2597 1392 -2596 ne
rect 1392 -2597 1393 -2596
tri 1393 -2597 1395 -2596 sw
tri 1401 -2597 1403 -2596 se
rect 395 -2600 396 -2599
tri 396 -2600 398 -2599 sw
tri 398 -2600 400 -2599 se
tri 395 -2602 396 -2600 ne
rect -604 -2605 -603 -2604
tri -603 -2605 -602 -2604 nw
tri -602 -2605 -601 -2604 ne
rect -601 -2605 -600 -2604
tri -600 -2605 -597 -2602 sw
tri 393 -2605 396 -2602 se
rect 396 -2604 400 -2600
tri 400 -2602 403 -2599 nw
tri 1392 -2600 1395 -2597 ne
tri 1395 -2599 1396 -2597 sw
tri 1400 -2599 1401 -2597 se
rect 1401 -2599 1403 -2597
tri 1403 -2599 1406 -2596 nw
tri 2390 -2596 2392 -2594 se
tri 2392 -2596 2393 -2594 sw
tri 2403 -2596 2404 -2594 se
tri 2404 -2596 2406 -2594 sw
tri 2390 -2597 2392 -2596 ne
rect 2392 -2597 2393 -2596
tri 2393 -2597 2395 -2596 sw
tri 2401 -2597 2403 -2596 se
rect 1395 -2600 1396 -2599
tri 1396 -2600 1398 -2599 sw
tri 1398 -2600 1400 -2599 se
tri 1395 -2602 1396 -2600 ne
rect 396 -2605 397 -2604
tri 397 -2605 398 -2604 nw
tri 398 -2605 399 -2604 ne
rect 399 -2605 400 -2604
tri 400 -2605 403 -2602 sw
tri 1393 -2605 1396 -2602 se
rect 1396 -2604 1400 -2600
tri 1400 -2602 1403 -2599 nw
tri 2392 -2600 2395 -2597 ne
tri 2395 -2599 2396 -2597 sw
tri 2400 -2599 2401 -2597 se
rect 2401 -2599 2403 -2597
tri 2403 -2599 2406 -2596 nw
tri 3390 -2596 3392 -2594 se
tri 3392 -2596 3393 -2594 sw
tri 3403 -2596 3404 -2594 se
tri 3404 -2596 3406 -2594 sw
tri 3390 -2597 3392 -2596 ne
rect 3392 -2597 3393 -2596
tri 3393 -2597 3395 -2596 sw
tri 3401 -2597 3403 -2596 se
rect 2395 -2600 2396 -2599
tri 2396 -2600 2398 -2599 sw
tri 2398 -2600 2400 -2599 se
tri 2395 -2602 2396 -2600 ne
rect 1396 -2605 1397 -2604
tri 1397 -2605 1398 -2604 nw
tri 1398 -2605 1399 -2604 ne
rect 1399 -2605 1400 -2604
tri 1400 -2605 1403 -2602 sw
tri 2393 -2605 2396 -2602 se
rect 2396 -2604 2400 -2600
tri 2400 -2602 2403 -2599 nw
tri 3392 -2600 3395 -2597 ne
tri 3395 -2599 3396 -2597 sw
tri 3400 -2599 3401 -2597 se
rect 3401 -2599 3403 -2597
tri 3403 -2599 3406 -2596 nw
rect 3395 -2600 3396 -2599
tri 3396 -2600 3398 -2599 sw
tri 3398 -2600 3400 -2599 se
tri 3395 -2602 3396 -2600 ne
rect 2396 -2605 2397 -2604
tri 2397 -2605 2398 -2604 nw
tri 2398 -2605 2399 -2604 ne
rect 2399 -2605 2400 -2604
tri 2400 -2605 2403 -2602 sw
tri 3393 -2605 3396 -2602 se
rect 3396 -2604 3400 -2600
tri 3400 -2602 3403 -2599 nw
rect 3396 -2605 3397 -2604
tri 3397 -2605 3398 -2604 nw
tri 3398 -2605 3399 -2604 ne
rect 3399 -2605 3400 -2604
tri 3400 -2605 3403 -2602 sw
tri -610 -2608 -607 -2605 se
tri -607 -2608 -604 -2605 nw
tri -600 -2608 -597 -2605 ne
tri -597 -2608 -594 -2605 sw
tri -610 -2610 -608 -2608 ne
tri -608 -2610 -607 -2608 nw
tri -597 -2610 -596 -2608 ne
tri -596 -2610 -594 -2608 nw
tri 390 -2608 393 -2605 se
tri 393 -2608 396 -2605 nw
tri 400 -2608 403 -2605 ne
tri 403 -2608 406 -2605 sw
tri 390 -2610 392 -2608 ne
tri 392 -2610 393 -2608 nw
tri 403 -2610 404 -2608 ne
tri 404 -2610 406 -2608 nw
tri 1390 -2608 1393 -2605 se
tri 1393 -2608 1396 -2605 nw
tri 1400 -2608 1403 -2605 ne
tri 1403 -2608 1406 -2605 sw
tri 1390 -2610 1392 -2608 ne
tri 1392 -2610 1393 -2608 nw
tri 1403 -2610 1404 -2608 ne
tri 1404 -2610 1406 -2608 nw
tri 2390 -2608 2393 -2605 se
tri 2393 -2608 2396 -2605 nw
tri 2400 -2608 2403 -2605 ne
tri 2403 -2608 2406 -2605 sw
tri 2390 -2610 2392 -2608 ne
tri 2392 -2610 2393 -2608 nw
tri 2403 -2610 2404 -2608 ne
tri 2404 -2610 2406 -2608 nw
tri 3390 -2608 3393 -2605 se
tri 3393 -2608 3396 -2605 nw
tri 3400 -2608 3403 -2605 ne
tri 3403 -2608 3406 -2605 sw
tri 3390 -2610 3392 -2608 ne
tri 3392 -2610 3393 -2608 nw
tri 3403 -2610 3404 -2608 ne
tri 3404 -2610 3406 -2608 nw
rect -534 -2670 -533 -2657
tri -533 -2670 -529 -2666 se
tri -470 -2670 -466 -2666 sw
rect -466 -2670 -465 -2657
rect -534 -2671 -465 -2670
rect -534 -2683 -533 -2671
tri -533 -2675 -529 -2671 ne
tri -470 -2675 -466 -2671 nw
rect -466 -2683 -465 -2671
rect -331 -2670 -330 -2657
tri -330 -2670 -326 -2666 se
tri -235 -2670 -231 -2666 sw
rect -231 -2670 -230 -2657
rect -331 -2671 -230 -2670
rect -331 -2683 -330 -2671
tri -330 -2675 -326 -2671 ne
tri -235 -2675 -231 -2671 nw
rect -231 -2683 -230 -2671
rect 466 -2670 467 -2657
tri 467 -2670 471 -2666 se
tri 530 -2670 534 -2666 sw
rect 534 -2670 535 -2657
rect 466 -2671 535 -2670
rect 466 -2683 467 -2671
tri 467 -2675 471 -2671 ne
tri 530 -2675 534 -2671 nw
rect 534 -2683 535 -2671
rect 669 -2670 670 -2657
tri 670 -2670 674 -2666 se
tri 765 -2670 769 -2666 sw
rect 769 -2670 770 -2657
rect 669 -2671 770 -2670
rect 669 -2683 670 -2671
tri 670 -2675 674 -2671 ne
tri 765 -2675 769 -2671 nw
rect 769 -2683 770 -2671
rect 1466 -2670 1467 -2657
tri 1467 -2670 1471 -2666 se
tri 1530 -2670 1534 -2666 sw
rect 1534 -2670 1535 -2657
rect 1466 -2671 1535 -2670
rect 1466 -2683 1467 -2671
tri 1467 -2675 1471 -2671 ne
tri 1530 -2675 1534 -2671 nw
rect 1534 -2683 1535 -2671
rect 1669 -2670 1670 -2657
tri 1670 -2670 1674 -2666 se
tri 1765 -2670 1769 -2666 sw
rect 1769 -2670 1770 -2657
rect 1669 -2671 1770 -2670
rect 1669 -2683 1670 -2671
tri 1670 -2675 1674 -2671 ne
tri 1765 -2675 1769 -2671 nw
rect 1769 -2683 1770 -2671
rect 2466 -2670 2467 -2657
tri 2467 -2670 2471 -2666 se
tri 2530 -2670 2534 -2666 sw
rect 2534 -2670 2535 -2657
rect 2466 -2671 2535 -2670
rect 2466 -2683 2467 -2671
tri 2467 -2675 2471 -2671 ne
tri 2530 -2675 2534 -2671 nw
rect 2534 -2683 2535 -2671
rect 2669 -2670 2670 -2657
tri 2670 -2670 2674 -2666 se
tri 2765 -2670 2769 -2666 sw
rect 2769 -2670 2770 -2657
rect 2669 -2671 2770 -2670
rect 2669 -2683 2670 -2671
tri 2670 -2675 2674 -2671 ne
tri 2765 -2675 2769 -2671 nw
rect 2769 -2683 2770 -2671
rect 3466 -2670 3467 -2657
tri 3467 -2670 3471 -2666 se
tri 3530 -2670 3534 -2666 sw
rect 3534 -2670 3535 -2657
rect 3466 -2671 3535 -2670
rect 3466 -2683 3467 -2671
tri 3467 -2675 3471 -2671 ne
tri 3530 -2675 3534 -2671 nw
rect 3534 -2683 3535 -2671
rect 3669 -2670 3670 -2657
tri 3670 -2670 3674 -2666 se
tri 3765 -2670 3769 -2666 sw
rect 3769 -2670 3770 -2657
rect 3669 -2671 3770 -2670
rect 3669 -2683 3670 -2671
tri 3670 -2675 3674 -2671 ne
tri 3765 -2675 3769 -2671 nw
rect 3769 -2683 3770 -2671
rect -811 -2824 -810 -2811
tri -810 -2824 -806 -2820 se
tri -398 -2824 -394 -2820 sw
rect -394 -2824 -393 -2811
rect -811 -2825 -623 -2824
rect -581 -2825 -393 -2824
rect -811 -2837 -810 -2825
tri -810 -2829 -806 -2825 ne
tri -398 -2829 -394 -2825 nw
rect -394 -2837 -393 -2825
rect 189 -2824 190 -2811
tri 190 -2824 194 -2820 se
tri 602 -2824 606 -2820 sw
rect 606 -2824 607 -2811
rect 189 -2825 377 -2824
rect 419 -2825 607 -2824
rect 189 -2837 190 -2825
tri 190 -2829 194 -2825 ne
tri 602 -2829 606 -2825 nw
rect 606 -2837 607 -2825
rect 1189 -2824 1190 -2811
tri 1190 -2824 1194 -2820 se
tri 1602 -2824 1606 -2820 sw
rect 1606 -2824 1607 -2811
rect 1189 -2825 1377 -2824
rect 1419 -2825 1607 -2824
rect 1189 -2837 1190 -2825
tri 1190 -2829 1194 -2825 ne
tri 1602 -2829 1606 -2825 nw
rect 1606 -2837 1607 -2825
rect 2189 -2824 2190 -2811
tri 2190 -2824 2194 -2820 se
tri 2602 -2824 2606 -2820 sw
rect 2606 -2824 2607 -2811
rect 2189 -2825 2377 -2824
rect 2419 -2825 2607 -2824
rect 2189 -2837 2190 -2825
tri 2190 -2829 2194 -2825 ne
tri 2602 -2829 2606 -2825 nw
rect 2606 -2837 2607 -2825
rect 3189 -2824 3190 -2811
tri 3190 -2824 3194 -2820 se
tri 3602 -2824 3606 -2820 sw
rect 3606 -2824 3607 -2811
rect 3189 -2825 3377 -2824
rect 3419 -2825 3607 -2824
rect 3189 -2837 3190 -2825
tri 3190 -2829 3194 -2825 ne
tri 3602 -2829 3606 -2825 nw
rect 3606 -2837 3607 -2825
rect -638 -2864 -637 -2851
tri -637 -2864 -633 -2860 se
tri -571 -2864 -567 -2860 sw
rect -567 -2864 -566 -2851
rect -638 -2865 -566 -2864
rect -638 -2877 -637 -2865
tri -637 -2869 -633 -2865 ne
tri -571 -2869 -567 -2865 nw
rect -567 -2877 -566 -2865
rect 362 -2864 363 -2851
tri 363 -2864 367 -2860 se
tri 429 -2864 433 -2860 sw
rect 433 -2864 434 -2851
rect 362 -2865 434 -2864
rect 362 -2877 363 -2865
tri 363 -2869 367 -2865 ne
tri 429 -2869 433 -2865 nw
rect 433 -2877 434 -2865
rect 1362 -2864 1363 -2851
tri 1363 -2864 1367 -2860 se
tri 1429 -2864 1433 -2860 sw
rect 1433 -2864 1434 -2851
rect 1362 -2865 1434 -2864
rect 1362 -2877 1363 -2865
tri 1363 -2869 1367 -2865 ne
tri 1429 -2869 1433 -2865 nw
rect 1433 -2877 1434 -2865
rect 2362 -2864 2363 -2851
tri 2363 -2864 2367 -2860 se
tri 2429 -2864 2433 -2860 sw
rect 2433 -2864 2434 -2851
rect 2362 -2865 2434 -2864
rect 2362 -2877 2363 -2865
tri 2363 -2869 2367 -2865 ne
tri 2429 -2869 2433 -2865 nw
rect 2433 -2877 2434 -2865
rect 3362 -2864 3363 -2851
tri 3363 -2864 3367 -2860 se
tri 3429 -2864 3433 -2860 sw
rect 3433 -2864 3434 -2851
rect 3362 -2865 3434 -2864
rect 3362 -2877 3363 -2865
tri 3363 -2869 3367 -2865 ne
tri 3429 -2869 3433 -2865 nw
rect 3433 -2877 3434 -2865
use sky130_fd_pr__pnp_05v5_W0p68L0p68  sky130_fd_pr__pnp_05v5_W0p68L0p68_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1620268331
transform 1 0 0 0 1 0
box 0 0 796 796
<< labels >>
flabel locali s 1375 378 1421 422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 1702 383 1743 409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 1556 384 1583 410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 1405 90 1405 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 1405 223 1405 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 1169 517 1169 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 1169 496 1169 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 1397 148 1397 148 0 FreeSans 100 0 0 0 0.360
flabel comment s 1398 784 1398 784 0 FreeSans 100 0 0 0 3.720
flabel comment s 1398 621 1398 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 1719 342 1719 342 0 FreeSans 100 0 0 0 0.505
flabel comment s 1638 545 1638 545 0 FreeSans 100 0 0 0 0.310
flabel comment s 1224 454 1224 454 0 FreeSans 100 0 0 0 0.360
flabel comment s 1500 342 1500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s 1398 177 1398 177 0 FreeSans 100 0 0 0 2.090
flabel comment s 1398 480 1398 480 0 FreeSans 100 0 0 0 0.068
flabel locali s 2375 378 2421 422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 2702 383 2743 409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 2556 384 2583 410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 2405 90 2405 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 2405 223 2405 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 2169 517 2169 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 2169 496 2169 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 2397 148 2397 148 0 FreeSans 100 0 0 0 0.360
flabel comment s 2398 784 2398 784 0 FreeSans 100 0 0 0 3.720
flabel comment s 2398 621 2398 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 2719 342 2719 342 0 FreeSans 100 0 0 0 0.505
flabel comment s 2638 545 2638 545 0 FreeSans 100 0 0 0 0.310
flabel comment s 2224 454 2224 454 0 FreeSans 100 0 0 0 0.360
flabel comment s 2500 342 2500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s 2398 177 2398 177 0 FreeSans 100 0 0 0 2.090
flabel comment s 2398 480 2398 480 0 FreeSans 100 0 0 0 0.068
flabel locali s 1375 -622 1421 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 1702 -617 1743 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 1556 -616 1583 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 1405 -910 1405 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 1405 -777 1405 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 1169 -483 1169 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 1169 -504 1169 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 1397 -852 1397 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s 1398 -216 1398 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s 1398 -379 1398 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 1719 -658 1719 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s 1638 -455 1638 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s 1224 -546 1224 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s 1500 -658 1500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s 1398 -823 1398 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s 1398 -520 1398 -520 0 FreeSans 100 0 0 0 0.068
flabel locali s 2375 -622 2421 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 2702 -617 2743 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 2556 -616 2583 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 2405 -910 2405 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 2405 -777 2405 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 2169 -483 2169 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 2169 -504 2169 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 2397 -852 2397 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s 2398 -216 2398 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s 2398 -379 2398 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 2719 -658 2719 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s 2638 -455 2638 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s 2224 -546 2224 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s 2500 -658 2500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s 2398 -823 2398 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s 2398 -520 2398 -520 0 FreeSans 100 0 0 0 0.068
flabel comment s 398 -520 398 -520 0 FreeSans 100 0 0 0 0.068
flabel comment s 398 -823 398 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s 500 -658 500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s 224 -546 224 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s 638 -455 638 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s 719 -658 719 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s 398 -379 398 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 398 -216 398 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s 397 -852 397 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s 169 -504 169 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 169 -483 169 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 405 -777 405 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 405 -910 405 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s 556 -616 583 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s 702 -617 743 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 375 -622 421 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 1375 -1622 1421 -1578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 1702 -1617 1743 -1591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 1556 -1616 1583 -1590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 1405 -1910 1405 -1910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 1405 -1777 1405 -1777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 1169 -1483 1169 -1483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 1169 -1504 1169 -1504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 1397 -1852 1397 -1852 0 FreeSans 100 0 0 0 0.360
flabel comment s 1398 -1216 1398 -1216 0 FreeSans 100 0 0 0 3.720
flabel comment s 1398 -1379 1398 -1379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 1719 -1658 1719 -1658 0 FreeSans 100 0 0 0 0.505
flabel comment s 1638 -1455 1638 -1455 0 FreeSans 100 0 0 0 0.310
flabel comment s 1224 -1546 1224 -1546 0 FreeSans 100 0 0 0 0.360
flabel comment s 1500 -1658 1500 -1658 0 FreeSans 100 0 0 0 0.345
flabel comment s 1398 -1823 1398 -1823 0 FreeSans 100 0 0 0 2.090
flabel comment s 1398 -1520 1398 -1520 0 FreeSans 100 0 0 0 0.068
flabel locali s 2375 -1622 2421 -1578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 2702 -1617 2743 -1591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 2556 -1616 2583 -1590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 2405 -1910 2405 -1910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 2405 -1777 2405 -1777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 2169 -1483 2169 -1483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 2169 -1504 2169 -1504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 2397 -1852 2397 -1852 0 FreeSans 100 0 0 0 0.360
flabel comment s 2398 -1216 2398 -1216 0 FreeSans 100 0 0 0 3.720
flabel comment s 2398 -1379 2398 -1379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 2719 -1658 2719 -1658 0 FreeSans 100 0 0 0 0.505
flabel comment s 2638 -1455 2638 -1455 0 FreeSans 100 0 0 0 0.310
flabel comment s 2224 -1546 2224 -1546 0 FreeSans 100 0 0 0 0.360
flabel comment s 2500 -1658 2500 -1658 0 FreeSans 100 0 0 0 0.345
flabel comment s 2398 -1823 2398 -1823 0 FreeSans 100 0 0 0 2.090
flabel comment s 2398 -1520 2398 -1520 0 FreeSans 100 0 0 0 0.068
flabel comment s 398 -1520 398 -1520 0 FreeSans 100 0 0 0 0.068
flabel comment s 398 -1823 398 -1823 0 FreeSans 100 0 0 0 2.090
flabel comment s 500 -1658 500 -1658 0 FreeSans 100 0 0 0 0.345
flabel comment s 224 -1546 224 -1546 0 FreeSans 100 0 0 0 0.360
flabel comment s 638 -1455 638 -1455 0 FreeSans 100 0 0 0 0.310
flabel comment s 719 -1658 719 -1658 0 FreeSans 100 0 0 0 0.505
flabel comment s 398 -1379 398 -1379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 398 -1216 398 -1216 0 FreeSans 100 0 0 0 3.720
flabel comment s 397 -1852 397 -1852 0 FreeSans 100 0 0 0 0.360
flabel comment s 169 -1504 169 -1504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 169 -1483 169 -1483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 405 -1777 405 -1777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 405 -1910 405 -1910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s 556 -1616 583 -1590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s 702 -1617 743 -1591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 375 -1622 421 -1578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -625 -1622 -579 -1578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -298 -1617 -257 -1591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -444 -1616 -417 -1590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s -595 -1910 -595 -1910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s -595 -1777 -595 -1777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -831 -1483 -831 -1483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -831 -1504 -831 -1504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -603 -1852 -603 -1852 0 FreeSans 100 0 0 0 0.360
flabel comment s -602 -1216 -602 -1216 0 FreeSans 100 0 0 0 3.720
flabel comment s -602 -1379 -602 -1379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -281 -1658 -281 -1658 0 FreeSans 100 0 0 0 0.505
flabel comment s -362 -1455 -362 -1455 0 FreeSans 100 0 0 0 0.310
flabel comment s -776 -1546 -776 -1546 0 FreeSans 100 0 0 0 0.360
flabel comment s -500 -1658 -500 -1658 0 FreeSans 100 0 0 0 0.345
flabel comment s -602 -1823 -602 -1823 0 FreeSans 100 0 0 0 2.090
flabel comment s -602 -1520 -602 -1520 0 FreeSans 100 0 0 0 0.068
flabel locali s 375 1378 421 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 702 1383 743 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 556 1384 583 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 405 1090 405 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 405 1223 405 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 169 1517 169 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 169 1496 169 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 397 1148 397 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s 398 1784 398 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s 398 1621 398 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 719 1342 719 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s 638 1545 638 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s 224 1454 224 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s 500 1342 500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s 398 1177 398 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s 398 1480 398 1480 0 FreeSans 100 0 0 0 0.068
flabel locali s 1375 1378 1421 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 1702 1383 1743 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 1556 1384 1583 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 1405 1090 1405 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 1405 1223 1405 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 1169 1517 1169 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 1169 1496 1169 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 1397 1148 1397 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s 1398 1784 1398 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s 1398 1621 1398 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 1719 1342 1719 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s 1638 1545 1638 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s 1224 1454 1224 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s 1500 1342 1500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s 1398 1177 1398 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s 1398 1480 1398 1480 0 FreeSans 100 0 0 0 0.068
flabel locali s 2375 1378 2421 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 2702 1383 2743 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 2556 1384 2583 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 2405 1090 2405 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 2405 1223 2405 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 2169 1517 2169 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 2169 1496 2169 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 2397 1148 2397 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s 2398 1784 2398 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s 2398 1621 2398 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 2719 1342 2719 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s 2638 1545 2638 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s 2224 1454 2224 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s 2500 1342 2500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s 2398 1177 2398 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s 2398 1480 2398 1480 0 FreeSans 100 0 0 0 0.068
flabel locali s 3375 1378 3421 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 3702 1383 3743 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 3556 1384 3583 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 3405 1090 3405 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 3405 1223 3405 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 3169 1517 3169 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 3169 1496 3169 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 3397 1148 3397 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s 3398 1784 3398 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s 3398 1621 3398 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 3719 1342 3719 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s 3638 1545 3638 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s 3224 1454 3224 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s 3500 1342 3500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s 3398 1177 3398 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s 3398 1480 3398 1480 0 FreeSans 100 0 0 0 0.068
flabel locali s 3375 378 3421 422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 3702 383 3743 409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 3556 384 3583 410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 3405 90 3405 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 3405 223 3405 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 3169 517 3169 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 3169 496 3169 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 3397 148 3397 148 0 FreeSans 100 0 0 0 0.360
flabel comment s 3398 784 3398 784 0 FreeSans 100 0 0 0 3.720
flabel comment s 3398 621 3398 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 3719 342 3719 342 0 FreeSans 100 0 0 0 0.505
flabel comment s 3638 545 3638 545 0 FreeSans 100 0 0 0 0.310
flabel comment s 3224 454 3224 454 0 FreeSans 100 0 0 0 0.360
flabel comment s 3500 342 3500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s 3398 177 3398 177 0 FreeSans 100 0 0 0 2.090
flabel comment s 3398 480 3398 480 0 FreeSans 100 0 0 0 0.068
flabel locali s 3375 -622 3421 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 3702 -617 3743 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 3556 -616 3583 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 3405 -910 3405 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 3405 -777 3405 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 3169 -483 3169 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 3169 -504 3169 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 3397 -852 3397 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s 3398 -216 3398 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s 3398 -379 3398 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 3719 -658 3719 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s 3638 -455 3638 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s 3224 -546 3224 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s 3500 -658 3500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s 3398 -823 3398 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s 3398 -520 3398 -520 0 FreeSans 100 0 0 0 0.068
flabel locali s 3375 -1622 3421 -1578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 3702 -1617 3743 -1591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 3556 -1616 3583 -1590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 3405 -1910 3405 -1910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 3405 -1777 3405 -1777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 3169 -1483 3169 -1483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 3169 -1504 3169 -1504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 3397 -1852 3397 -1852 0 FreeSans 100 0 0 0 0.360
flabel comment s 3398 -1216 3398 -1216 0 FreeSans 100 0 0 0 3.720
flabel comment s 3398 -1379 3398 -1379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 3719 -1658 3719 -1658 0 FreeSans 100 0 0 0 0.505
flabel comment s 3638 -1455 3638 -1455 0 FreeSans 100 0 0 0 0.310
flabel comment s 3224 -1546 3224 -1546 0 FreeSans 100 0 0 0 0.360
flabel comment s 3500 -1658 3500 -1658 0 FreeSans 100 0 0 0 0.345
flabel comment s 3398 -1823 3398 -1823 0 FreeSans 100 0 0 0 2.090
flabel comment s 3398 -1520 3398 -1520 0 FreeSans 100 0 0 0 0.068
flabel locali s 3375 -2622 3421 -2578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 3702 -2617 3743 -2591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 3556 -2616 3583 -2590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 3405 -2910 3405 -2910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 3405 -2777 3405 -2777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 3169 -2483 3169 -2483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 3169 -2504 3169 -2504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 3397 -2852 3397 -2852 0 FreeSans 100 0 0 0 0.360
flabel comment s 3398 -2216 3398 -2216 0 FreeSans 100 0 0 0 3.720
flabel comment s 3398 -2379 3398 -2379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 3719 -2658 3719 -2658 0 FreeSans 100 0 0 0 0.505
flabel comment s 3638 -2455 3638 -2455 0 FreeSans 100 0 0 0 0.310
flabel comment s 3224 -2546 3224 -2546 0 FreeSans 100 0 0 0 0.360
flabel comment s 3500 -2658 3500 -2658 0 FreeSans 100 0 0 0 0.345
flabel comment s 3398 -2823 3398 -2823 0 FreeSans 100 0 0 0 2.090
flabel comment s 3398 -2520 3398 -2520 0 FreeSans 100 0 0 0 0.068
flabel locali s 2375 -2622 2421 -2578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 2702 -2617 2743 -2591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 2556 -2616 2583 -2590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 2405 -2910 2405 -2910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 2405 -2777 2405 -2777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 2169 -2483 2169 -2483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 2169 -2504 2169 -2504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 2397 -2852 2397 -2852 0 FreeSans 100 0 0 0 0.360
flabel comment s 2398 -2216 2398 -2216 0 FreeSans 100 0 0 0 3.720
flabel comment s 2398 -2379 2398 -2379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 2719 -2658 2719 -2658 0 FreeSans 100 0 0 0 0.505
flabel comment s 2638 -2455 2638 -2455 0 FreeSans 100 0 0 0 0.310
flabel comment s 2224 -2546 2224 -2546 0 FreeSans 100 0 0 0 0.360
flabel comment s 2500 -2658 2500 -2658 0 FreeSans 100 0 0 0 0.345
flabel comment s 2398 -2823 2398 -2823 0 FreeSans 100 0 0 0 2.090
flabel comment s 2398 -2520 2398 -2520 0 FreeSans 100 0 0 0 0.068
flabel locali s 1375 -2622 1421 -2578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 1702 -2617 1743 -2591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 1556 -2616 1583 -2590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 1405 -2910 1405 -2910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 1405 -2777 1405 -2777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 1169 -2483 1169 -2483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 1169 -2504 1169 -2504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 1397 -2852 1397 -2852 0 FreeSans 100 0 0 0 0.360
flabel comment s 1398 -2216 1398 -2216 0 FreeSans 100 0 0 0 3.720
flabel comment s 1398 -2379 1398 -2379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 1719 -2658 1719 -2658 0 FreeSans 100 0 0 0 0.505
flabel comment s 1638 -2455 1638 -2455 0 FreeSans 100 0 0 0 0.310
flabel comment s 1224 -2546 1224 -2546 0 FreeSans 100 0 0 0 0.360
flabel comment s 1500 -2658 1500 -2658 0 FreeSans 100 0 0 0 0.345
flabel comment s 1398 -2823 1398 -2823 0 FreeSans 100 0 0 0 2.090
flabel comment s 1398 -2520 1398 -2520 0 FreeSans 100 0 0 0 0.068
flabel locali s 375 -2622 421 -2578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 702 -2617 743 -2591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 556 -2616 583 -2590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 405 -2910 405 -2910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 405 -2777 405 -2777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 169 -2483 169 -2483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 169 -2504 169 -2504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 397 -2852 397 -2852 0 FreeSans 100 0 0 0 0.360
flabel comment s 398 -2216 398 -2216 0 FreeSans 100 0 0 0 3.720
flabel comment s 398 -2379 398 -2379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 719 -2658 719 -2658 0 FreeSans 100 0 0 0 0.505
flabel comment s 638 -2455 638 -2455 0 FreeSans 100 0 0 0 0.310
flabel comment s 224 -2546 224 -2546 0 FreeSans 100 0 0 0 0.360
flabel comment s 500 -2658 500 -2658 0 FreeSans 100 0 0 0 0.345
flabel comment s 398 -2823 398 -2823 0 FreeSans 100 0 0 0 2.090
flabel comment s 398 -2520 398 -2520 0 FreeSans 100 0 0 0 0.068
flabel locali s -625 -2622 -579 -2578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -298 -2617 -257 -2591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -444 -2616 -417 -2590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s -595 -2910 -595 -2910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s -595 -2777 -595 -2777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -831 -2483 -831 -2483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -831 -2504 -831 -2504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -603 -2852 -603 -2852 0 FreeSans 100 0 0 0 0.360
flabel comment s -602 -2216 -602 -2216 0 FreeSans 100 0 0 0 3.720
flabel comment s -602 -2379 -602 -2379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -281 -2658 -281 -2658 0 FreeSans 100 0 0 0 0.505
flabel comment s -362 -2455 -362 -2455 0 FreeSans 100 0 0 0 0.310
flabel comment s -776 -2546 -776 -2546 0 FreeSans 100 0 0 0 0.360
flabel comment s -500 -2658 -500 -2658 0 FreeSans 100 0 0 0 0.345
flabel comment s -602 -2823 -602 -2823 0 FreeSans 100 0 0 0 2.090
flabel comment s -602 -2520 -602 -2520 0 FreeSans 100 0 0 0 0.068
flabel comment s -602 1480 -602 1480 0 FreeSans 100 0 0 0 0.068
flabel comment s -602 1177 -602 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s -500 1342 -500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s -776 1454 -776 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s -362 1545 -362 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s -281 1342 -281 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s -602 1621 -602 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -602 1784 -602 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s -603 1148 -603 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s -831 1496 -831 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -831 1517 -831 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -595 1223 -595 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -595 1090 -595 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -444 1384 -417 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -298 1383 -257 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -625 1378 -579 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel comment s -602 -520 -602 -520 0 FreeSans 100 0 0 0 0.068
flabel comment s -602 -823 -602 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s -500 -658 -500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s -776 -546 -776 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s -362 -455 -362 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s -281 -658 -281 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s -602 -379 -602 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -602 -216 -602 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s -603 -852 -603 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s -831 -504 -831 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -831 -483 -831 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -595 -777 -595 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -595 -910 -595 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -444 -616 -417 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -298 -617 -257 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -625 -622 -579 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel comment s -602 480 -602 480 0 FreeSans 100 0 0 0 0.068
flabel comment s -602 177 -602 177 0 FreeSans 100 0 0 0 2.090
flabel comment s -500 342 -500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s -776 454 -776 454 0 FreeSans 100 0 0 0 0.360
flabel comment s -362 545 -362 545 0 FreeSans 100 0 0 0 0.310
flabel comment s -281 342 -281 342 0 FreeSans 100 0 0 0 0.505
flabel comment s -602 621 -602 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -602 784 -602 784 0 FreeSans 100 0 0 0 3.720
flabel comment s -603 148 -603 148 0 FreeSans 100 0 0 0 0.360
flabel comment s -831 496 -831 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -831 517 -831 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -595 223 -595 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -595 90 -595 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -444 384 -417 410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -298 383 -257 409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -625 378 -579 422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -1625 378 -1579 422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -1298 383 -1257 409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -1444 384 -1417 410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s -1595 90 -1595 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s -1595 223 -1595 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -1831 517 -1831 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -1831 496 -1831 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -1603 148 -1603 148 0 FreeSans 100 0 0 0 0.360
flabel comment s -1602 784 -1602 784 0 FreeSans 100 0 0 0 3.720
flabel comment s -1602 621 -1602 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -1281 342 -1281 342 0 FreeSans 100 0 0 0 0.505
flabel comment s -1362 545 -1362 545 0 FreeSans 100 0 0 0 0.310
flabel comment s -1776 454 -1776 454 0 FreeSans 100 0 0 0 0.360
flabel comment s -1500 342 -1500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s -1602 177 -1602 177 0 FreeSans 100 0 0 0 2.090
flabel comment s -1602 480 -1602 480 0 FreeSans 100 0 0 0 0.068
flabel locali s -1625 -622 -1579 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -1298 -617 -1257 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -1444 -616 -1417 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s -1595 -910 -1595 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s -1595 -777 -1595 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -1831 -483 -1831 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -1831 -504 -1831 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -1603 -852 -1603 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s -1602 -216 -1602 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s -1602 -379 -1602 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -1281 -658 -1281 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s -1362 -455 -1362 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s -1776 -546 -1776 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s -1500 -658 -1500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s -1602 -823 -1602 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s -1602 -520 -1602 -520 0 FreeSans 100 0 0 0 0.068
flabel comment s -2602 -520 -2602 -520 0 FreeSans 100 0 0 0 0.068
flabel comment s -2602 -823 -2602 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s -2500 -658 -2500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s -2776 -546 -2776 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s -2362 -455 -2362 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s -2281 -658 -2281 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s -2602 -379 -2602 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -2602 -216 -2602 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s -2603 -852 -2603 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s -2831 -504 -2831 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -2831 -483 -2831 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -2595 -777 -2595 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -2595 -910 -2595 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -2444 -616 -2417 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -2298 -617 -2257 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -2625 -622 -2579 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -2625 1378 -2579 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -2298 1383 -2257 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -2444 1384 -2417 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s -2595 1090 -2595 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s -2595 1223 -2595 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -2831 1517 -2831 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -2831 1496 -2831 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -2603 1148 -2603 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s -2602 1784 -2602 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s -2602 1621 -2602 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -2281 1342 -2281 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s -2362 1545 -2362 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s -2776 1454 -2776 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s -2500 1342 -2500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s -2602 1177 -2602 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s -2602 1480 -2602 1480 0 FreeSans 100 0 0 0 0.068
flabel locali s -1625 1378 -1579 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s -1298 1383 -1257 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -1444 1384 -1417 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s -1595 1090 -1595 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s -1595 1223 -1595 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -1831 1517 -1831 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -1831 1496 -1831 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -1603 1148 -1603 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s -1602 1784 -1602 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s -1602 1621 -1602 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -1281 1342 -1281 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s -1362 1545 -1362 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s -1776 1454 -1776 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s -1500 1342 -1500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s -1602 1177 -1602 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s -1602 1480 -1602 1480 0 FreeSans 100 0 0 0 0.068
flabel comment s -3602 1480 -3602 1480 0 FreeSans 100 0 0 0 0.068
flabel comment s -3602 1177 -3602 1177 0 FreeSans 100 0 0 0 2.090
flabel comment s -3500 1342 -3500 1342 0 FreeSans 100 0 0 0 0.345
flabel comment s -3776 1454 -3776 1454 0 FreeSans 100 0 0 0 0.360
flabel comment s -3362 1545 -3362 1545 0 FreeSans 100 0 0 0 0.310
flabel comment s -3281 1342 -3281 1342 0 FreeSans 100 0 0 0 0.505
flabel comment s -3602 1621 -3602 1621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -3602 1784 -3602 1784 0 FreeSans 100 0 0 0 3.720
flabel comment s -3603 1148 -3603 1148 0 FreeSans 100 0 0 0 0.360
flabel comment s -3831 1496 -3831 1496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -3831 1517 -3831 1517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -3595 1223 -3595 1223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -3595 1090 -3595 1090 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -3444 1384 -3417 1410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -3298 1383 -3257 1409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -3625 1378 -3579 1422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel comment s -3602 -520 -3602 -520 0 FreeSans 100 0 0 0 0.068
flabel comment s -3602 -823 -3602 -823 0 FreeSans 100 0 0 0 2.090
flabel comment s -3500 -658 -3500 -658 0 FreeSans 100 0 0 0 0.345
flabel comment s -3776 -546 -3776 -546 0 FreeSans 100 0 0 0 0.360
flabel comment s -3362 -455 -3362 -455 0 FreeSans 100 0 0 0 0.310
flabel comment s -3281 -658 -3281 -658 0 FreeSans 100 0 0 0 0.505
flabel comment s -3602 -379 -3602 -379 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -3602 -216 -3602 -216 0 FreeSans 100 0 0 0 3.720
flabel comment s -3603 -852 -3603 -852 0 FreeSans 100 0 0 0 0.360
flabel comment s -3831 -504 -3831 -504 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -3831 -483 -3831 -483 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -3595 -777 -3595 -777 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -3595 -910 -3595 -910 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -3444 -616 -3417 -590 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -3298 -617 -3257 -591 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -3625 -622 -3579 -578 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel comment s -3602 480 -3602 480 0 FreeSans 100 0 0 0 0.068
flabel comment s -3602 177 -3602 177 0 FreeSans 100 0 0 0 2.090
flabel comment s -3500 342 -3500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s -3776 454 -3776 454 0 FreeSans 100 0 0 0 0.360
flabel comment s -3362 545 -3362 545 0 FreeSans 100 0 0 0 0.310
flabel comment s -3281 342 -3281 342 0 FreeSans 100 0 0 0 0.505
flabel comment s -3602 621 -3602 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -3602 784 -3602 784 0 FreeSans 100 0 0 0 3.720
flabel comment s -3603 148 -3603 148 0 FreeSans 100 0 0 0 0.360
flabel comment s -3831 496 -3831 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -3831 517 -3831 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -3595 223 -3595 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -3595 90 -3595 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -3444 384 -3417 410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -3298 383 -3257 409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -3625 378 -3579 422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel comment s -2602 480 -2602 480 0 FreeSans 100 0 0 0 0.068
flabel comment s -2602 177 -2602 177 0 FreeSans 100 0 0 0 2.090
flabel comment s -2500 342 -2500 342 0 FreeSans 100 0 0 0 0.345
flabel comment s -2776 454 -2776 454 0 FreeSans 100 0 0 0 0.360
flabel comment s -2362 545 -2362 545 0 FreeSans 100 0 0 0 0.310
flabel comment s -2281 342 -2281 342 0 FreeSans 100 0 0 0 0.505
flabel comment s -2602 621 -2602 621 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s -2602 784 -2602 784 0 FreeSans 100 0 0 0 3.720
flabel comment s -2603 148 -2603 148 0 FreeSans 100 0 0 0 0.360
flabel comment s -2831 496 -2831 496 0 FreeSans 100 0 0 0 adj. sides
flabel comment s -2831 517 -2831 517 0 FreeSans 100 0 0 0 0.12 min
flabel comment s -2595 223 -2595 223 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s -2595 90 -2595 90 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel locali s -2444 384 -2417 410 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel locali s -2298 383 -2257 409 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s -2625 378 -2579 422 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
<< end >>
