magic
tech sky130A
timestamp 1620687492
<< metal3 >>
rect -115 -15 415 515
<< mimcap >>
rect -100 295 400 500
rect -100 205 105 295
rect 195 205 400 295
rect -100 0 400 205
<< mimcapcontact >>
rect 105 205 195 295
<< metal4 >>
rect 100 295 200 300
rect 100 205 105 295
rect 195 205 200 295
rect 100 200 200 205
<< labels >>
rlabel metal3 415 40 415 40 3 2
rlabel metal4 200 245 200 245 3 1
<< end >>
