magic
tech sky130A
timestamp 1620604094
<< nwell >>
rect -90 1125 5 1365
rect 2645 1125 2680 1365
rect -90 465 5 705
rect 2645 465 2685 705
<< poly >>
rect 120 1490 2370 1505
rect -75 1455 -35 1465
rect -75 1435 -65 1455
rect -45 1435 -35 1455
rect -75 1425 -35 1435
rect -65 -20 -45 1425
rect 120 1360 135 1490
rect 1315 1390 1355 1400
rect 1315 1370 1325 1390
rect 1345 1370 1355 1390
rect 1315 1360 1355 1370
rect 2355 1360 2370 1490
rect 2605 1455 2645 1465
rect 2605 1435 2615 1455
rect 2635 1435 2645 1455
rect 2605 1425 2645 1435
rect 2605 1410 2665 1425
rect 1175 750 1355 765
rect 1340 740 1355 750
rect 1340 725 1525 740
rect 1340 700 1355 725
rect 1315 120 1355 130
rect 1180 95 1220 105
rect 1180 75 1190 95
rect 1210 75 1220 95
rect 1315 100 1325 120
rect 1345 100 1355 120
rect 1315 90 1355 100
rect 1180 65 1220 75
rect -75 -30 -35 -20
rect -75 -50 -65 -30
rect -45 -50 -35 -30
rect -75 -60 -35 -50
rect 1205 -65 1220 65
rect 1325 20 1345 90
rect 1315 10 1355 20
rect 1315 -10 1325 10
rect 1345 -10 1355 10
rect 1315 -20 1355 -10
rect 1545 0 1560 175
rect 1545 -10 1585 0
rect 1545 -30 1555 -10
rect 1575 -30 1585 -10
rect 1545 -40 1585 -30
rect 2650 -65 2665 1410
rect 1205 -80 2665 -65
<< polycont >>
rect -65 1435 -45 1455
rect 1325 1370 1345 1390
rect 2615 1435 2635 1455
rect 1190 75 1210 95
rect 1325 100 1345 120
rect -65 -50 -45 -30
rect 1325 -10 1345 10
rect 1555 -30 1575 -10
<< locali >>
rect -75 1455 -35 1465
rect -75 1445 -65 1455
rect -90 1435 -65 1445
rect -45 1445 -35 1455
rect 2605 1455 2645 1465
rect -45 1435 25 1445
rect -90 1425 25 1435
rect 2605 1435 2615 1455
rect 2635 1435 2645 1455
rect 2605 1425 2645 1435
rect -90 1380 25 1400
rect 1220 1390 1355 1400
rect 1220 1380 1325 1390
rect 1315 1370 1325 1380
rect 1345 1370 1355 1390
rect 1315 1360 1355 1370
rect 1380 1380 1440 1400
rect 2645 1380 2680 1400
rect 1380 1340 1400 1380
rect -90 835 45 855
rect 1520 720 1525 740
rect 1380 130 1400 185
rect 1315 120 1400 130
rect 1180 95 1220 105
rect -90 65 15 85
rect 1180 75 1190 95
rect 1210 75 1220 95
rect 1315 100 1325 120
rect 1345 110 1400 120
rect 1345 100 1355 110
rect 1315 90 1355 100
rect 1180 65 1220 75
rect 1375 65 1430 85
rect 2645 65 2680 85
rect 1375 60 1395 65
rect 1240 40 1395 60
rect 1240 -20 1260 40
rect 2645 20 2680 40
rect -75 -30 1260 -20
rect -75 -50 -65 -30
rect -45 -40 1260 -30
rect 1315 10 1355 20
rect 1315 -10 1325 10
rect 1345 -10 1355 10
rect -45 -50 -35 -40
rect -75 -60 -35 -50
rect 1315 -90 1355 -10
rect 1545 -10 1585 0
rect 1545 -30 1555 -10
rect 1575 -20 1585 -10
rect 1575 -30 2680 -20
rect 1545 -40 2680 -30
<< metal1 >>
rect -90 1150 30 1340
rect 2645 1150 2680 1340
rect -90 895 15 1085
rect 2645 895 2685 1085
rect -90 490 5 680
rect 2645 490 2685 680
rect -90 235 0 425
rect 2645 235 2685 425
use dff  dff_1
timestamp 1620594849
transform 1 0 1430 0 1 70
box -5 -70 1215 1395
use inverter  inverter_1
timestamp 1620435323
transform 1 0 1340 0 1 755
box -120 80 85 610
use inverter  inverter_0
timestamp 1620435323
transform 1 0 1340 0 1 95
box -120 80 85 610
use dff  dff_0
timestamp 1620594849
transform 1 0 5 0 1 70
box -5 -70 1215 1395
<< labels >>
rlabel locali 0 845 0 845 7 D
rlabel locali -90 1435 -90 1435 7 preset
rlabel locali -90 1390 -90 1390 7 clk
rlabel locali -90 845 -90 845 7 D
rlabel locali -90 75 -90 75 7 clear
rlabel metal1 -90 1245 -90 1245 7 VDD
rlabel metal1 -90 985 -90 985 7 GND
rlabel locali 2680 -30 2680 -30 3 Qout
rlabel locali 1335 -90 1335 -90 5 Qnout
<< end >>
