magic
tech sky130A
timestamp 1620704963
<< poly >>
rect -100 2600 20 2615
rect -100 -335 -85 2600
rect -10 -335 35 -325
rect -100 -350 0 -335
rect -10 -355 0 -350
rect 25 -355 35 -335
rect -10 -365 35 -355
<< polycont >>
rect 0 -355 25 -335
<< locali >>
rect 2875 -45 2920 595
rect 725 -65 2920 -45
rect -10 -335 35 -325
rect -10 -355 0 -335
rect 25 -355 35 -335
rect -10 -415 35 -355
rect 685 -415 725 -395
rect -10 -445 725 -415
rect 2875 -425 2920 -65
rect 2815 -445 2920 -425
rect 2815 -515 2835 -445
rect 2900 -515 2920 -445
rect 2815 -535 2920 -515
<< viali >>
rect 0 -355 25 -335
rect 2835 -515 2900 -445
<< metal1 >>
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -10 -365 35 -360
rect 2825 -445 2910 -435
rect 2825 -515 2835 -445
rect 2900 -515 2910 -445
rect 2825 -525 2910 -515
<< via1 >>
rect -5 -335 30 -330
rect -5 -355 0 -335
rect 0 -355 25 -335
rect 25 -355 30 -335
rect -5 -360 30 -355
rect 2835 -515 2900 -445
<< metal2 >>
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -10 -365 35 -360
rect 2825 -445 2910 -435
rect 2825 -515 2835 -445
rect 2900 -515 2910 -445
rect 2825 -525 2910 -515
<< via2 >>
rect -5 -360 30 -330
rect 2835 -515 2900 -445
<< metal3 >>
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -1525 -520 -1430 -390
rect -10 -520 35 -360
rect -1525 -555 35 -520
rect 2825 -445 2910 -435
rect 2825 -515 2835 -445
rect 2900 -515 2910 -445
rect 2825 -525 2910 -515
<< via3 >>
rect 2835 -515 2900 -445
<< metal4 >>
rect -1755 -425 -1630 -70
rect -1755 -445 2920 -425
rect -1755 -515 2835 -445
rect 2900 -515 2920 -445
rect -1755 -535 2920 -515
use switch  switch_0
timestamp 1620697026
transform 0 -1 1025 1 0 -290
box -110 20 245 625
use cap8to1  cap8to1_1
timestamp 1620703920
transform 1 0 -3915 0 1 1600
box 5 30 3785 1860
use cap8to1  cap8to1_0
timestamp 1620703920
transform 1 0 -3915 0 1 -430
box 5 30 3785 1860
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620692581
transform 1 0 255 0 1 -2315
box -255 2315 4445 5470
<< end >>
