magic
tech sky130A
timestamp 1620761386
<< poly >>
rect 7850 2910 7890 2920
rect 7850 2890 7860 2910
rect 7880 2895 7890 2910
rect 7880 2890 7910 2895
rect 7850 2880 7910 2890
rect -2145 2855 -2105 2865
rect -2145 2835 -2135 2855
rect -2115 2840 -2105 2855
rect 2865 2855 2905 2865
rect -2115 2835 -2085 2840
rect -2145 2825 -2085 2835
rect 2865 2835 2875 2855
rect 2895 2840 2905 2855
rect 2895 2835 2925 2840
rect 2865 2825 2925 2835
rect 7810 2160 7910 2170
rect 7810 2140 7820 2160
rect 7840 2155 7910 2160
rect 7840 2140 7850 2155
rect -2180 2130 -2140 2140
rect -2180 2110 -2170 2130
rect -2150 2115 -2140 2130
rect 2840 2130 2880 2140
rect 7810 2130 7850 2140
rect -2150 2110 -2070 2115
rect -2180 2100 -2070 2110
rect 2840 2110 2850 2130
rect 2870 2115 2880 2130
rect 2870 2110 2995 2115
rect 2840 2100 2995 2110
<< polycont >>
rect 7860 2890 7880 2910
rect -2135 2835 -2115 2855
rect 2875 2835 2895 2855
rect 7820 2140 7840 2160
rect -2170 2110 -2150 2130
rect 2850 2110 2870 2130
<< locali >>
rect 7850 3580 10890 3600
rect -2145 3495 895 3515
rect -2145 2865 -2125 3495
rect -2145 2855 -2105 2865
rect -2145 2835 -2135 2855
rect -2115 2835 -2105 2855
rect -2145 2825 -2105 2835
rect -2180 2130 -2140 2140
rect -2180 2110 -2170 2130
rect -2150 2110 -2140 2130
rect -2180 2100 -2140 2110
rect 875 795 895 3495
rect 2865 3495 5900 3515
rect 2865 2865 2885 3495
rect 2865 2855 2905 2865
rect 2865 2835 2875 2855
rect 2895 2835 2905 2855
rect 2865 2825 2905 2835
rect 2840 2130 2880 2140
rect 2840 2110 2850 2130
rect 2870 2110 2880 2130
rect 2840 210 2880 2110
rect 5880 795 5900 3495
rect 7850 2920 7870 3580
rect 7850 2910 7890 2920
rect 7850 2890 7860 2910
rect 7880 2890 7890 2910
rect 7850 2880 7890 2890
rect 7810 2160 7850 2170
rect 7810 2140 7820 2160
rect 7840 2140 7850 2160
rect 7810 2130 7850 2140
rect 2830 200 2880 210
rect 2830 175 2840 200
rect 2870 175 2880 200
rect 2830 165 2880 175
rect 7810 100 7830 2130
rect 10870 850 10890 3580
rect 4645 80 7830 100
rect 4645 -45 4695 80
<< viali >>
rect -2170 2110 -2150 2130
rect 2840 175 2870 200
<< metal1 >>
rect -2180 2130 -2140 2140
rect -2180 2110 -2170 2130
rect -2150 2110 -2140 2130
rect -2180 2100 -2140 2110
rect -2160 185 -2140 2100
rect 735 1030 1235 1040
rect 735 860 1165 1030
rect 1225 860 1235 1030
rect 735 850 1235 860
rect 5755 1030 6085 1040
rect 5755 860 5975 1030
rect 6075 860 6085 1030
rect 5755 850 6085 860
rect 750 600 3240 670
rect 195 575 3240 600
rect 195 495 3030 575
rect 5755 570 7990 655
rect 2830 200 2880 210
rect 2830 185 2840 200
rect -2160 175 2840 185
rect 2870 175 2880 200
rect -2160 165 2880 175
rect 2000 15 2080 165
rect 5285 -2360 8395 -2350
rect 5285 -2530 8120 -2360
rect 8380 -2530 8395 -2360
rect 5285 -2540 8395 -2530
rect 8595 -2625 9585 425
rect 5285 -2820 9585 -2625
<< via1 >>
rect 1165 860 1225 1030
rect 5975 860 6075 1030
rect 8120 -2530 8380 -2360
<< metal2 >>
rect 1155 1030 3035 1040
rect 1155 860 1165 1030
rect 1225 860 3035 1030
rect 1155 850 3035 860
rect 5965 1030 7985 1040
rect 5965 860 5975 1030
rect 6075 860 7985 1030
rect 5965 850 7985 860
rect 8105 -2360 8395 400
rect 8105 -2530 8120 -2360
rect 8380 -2530 8395 -2360
rect 8105 -2540 8395 -2530
use bandgap_thomas  bandgap_thomas_0
timestamp 1620761224
transform 1 0 -925 0 1 -3165
box 0 0 8070 3190
use selfbiasedcascode2stage  selfbiasedcascode2stage_1
timestamp 1620692581
transform 1 0 3170 0 1 -2090
box -255 2315 4445 5470
use selfbiasedcascode2stage  selfbiasedcascode2stage_2
timestamp 1620692581
transform 1 0 -1835 0 1 -2090
box -255 2315 4445 5470
use selfbiasedcascode2stage  selfbiasedcascode2stage_3
timestamp 1620692581
transform 1 0 8160 0 1 -2035
box -255 2315 4445 5470
<< end >>
