magic
tech sky130A
timestamp 1620759431
<< poly >>
rect 4355 2760 4580 2775
rect 5305 2750 5360 2760
rect 3520 2715 3570 2725
rect 3520 2690 3530 2715
rect 3560 2690 3570 2715
rect 5305 2715 5315 2750
rect 5350 2715 5360 2750
rect 5305 2705 5360 2715
rect 3520 2610 3570 2690
rect 3310 1910 3360 1920
rect 3310 1885 3320 1910
rect 3350 1890 3360 1910
rect 3350 1885 3380 1890
rect 3310 1875 3380 1885
<< polycont >>
rect 3530 2690 3560 2715
rect 5315 2715 5350 2750
rect 3320 1885 3350 1910
<< locali >>
rect 4640 3170 4690 3180
rect 4640 3145 4650 3170
rect 4680 3145 4690 3170
rect 4640 3080 4690 3145
rect 3310 1910 3360 2790
rect 3520 2715 3570 2805
rect 3520 2690 3530 2715
rect 3560 2690 3570 2715
rect 3520 2680 3570 2690
rect 4850 2720 4900 2805
rect 4850 2690 4860 2720
rect 4890 2690 4900 2720
rect 5305 2750 5360 2760
rect 5305 2715 5315 2750
rect 5350 2715 5360 2750
rect 5305 2705 5360 2715
rect 4850 2680 4900 2690
rect 3310 1885 3320 1910
rect 3350 1885 3360 1910
rect 3310 675 3360 1885
rect 3300 665 3360 675
rect 3300 635 3310 665
rect 3350 635 3360 665
rect 3300 625 3360 635
<< viali >>
rect 4650 3145 4680 3170
rect 3530 2690 3560 2715
rect 4860 2690 4890 2720
rect 5315 2715 5350 2750
rect 3310 635 3350 665
<< metal1 >>
rect 1405 3170 4690 3190
rect 1405 3150 4650 3170
rect 1405 2475 1495 3150
rect 4640 3145 4650 3150
rect 4680 3145 4690 3170
rect 4640 3135 4690 3145
rect 3320 2800 3350 3070
rect 4410 2790 4465 3080
rect 5305 2750 5360 2760
rect 2430 2715 3570 2725
rect 2430 2690 3530 2715
rect 3560 2690 3570 2715
rect 2430 2680 3570 2690
rect 4850 2720 4900 2730
rect 4850 2690 4860 2720
rect 4890 2690 4900 2720
rect 5305 2715 5315 2750
rect 5350 2715 5360 2750
rect 5305 2705 5360 2715
rect 4850 2680 4900 2690
rect 2160 2210 2240 2220
rect 2160 2165 2170 2210
rect 2230 2165 2240 2210
rect 2160 1900 2240 2165
rect 2430 1735 2475 2680
rect 5450 2640 5540 2800
rect 5370 2630 5540 2640
rect 5370 2595 5380 2630
rect 5530 2595 5540 2630
rect 5370 2585 5540 2595
rect 2160 1715 2475 1735
rect 2160 1400 2240 1715
rect 3300 665 3360 675
rect 3300 660 3310 665
rect 2045 635 3310 660
rect 3350 635 3360 665
rect 2045 625 3360 635
rect 2045 590 2155 625
<< via1 >>
rect 4860 2690 4890 2720
rect 5315 2715 5350 2750
rect 2170 2165 2230 2210
rect 5380 2595 5530 2630
<< metal2 >>
rect 5305 2750 5360 2760
rect 3265 2720 4900 2730
rect 3265 2690 4860 2720
rect 4890 2690 4900 2720
rect 5305 2715 5315 2750
rect 5350 2715 5360 2750
rect 5305 2705 5360 2715
rect 3265 2680 4900 2690
rect 3265 2220 3305 2680
rect 5370 2630 5540 2640
rect 5370 2595 5380 2630
rect 5530 2595 5540 2630
rect 5370 2505 5540 2595
rect 2160 2210 3305 2220
rect 2160 2165 2170 2210
rect 2230 2165 3305 2210
rect 2160 2155 3305 2165
<< via2 >>
rect 5315 2715 5350 2750
<< metal3 >>
rect 5305 2750 5845 2760
rect 5305 2715 5315 2750
rect 5350 2730 5845 2750
rect 5350 2715 5360 2730
rect 5305 2705 5360 2715
use bandgap_pnp_thomas  bandgap_pnp_thomas_0
timestamp 1620712167
transform 1 0 2000 0 1 2240
box -2000 -2240 1155 898
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620692581
transform 1 0 3625 0 1 -2315
box -255 2315 4445 5470
use bandgap_current_mirror  bandgap_current_mirror_0
timestamp 1620755988
transform 1 0 3240 0 1 2730
box -135 30 1195 390
use bandgap_current_mirror  bandgap_current_mirror_1
timestamp 1620755988
transform 1 0 4570 0 1 2730
box -135 30 1195 390
<< end >>
