magic
tech sky130A
timestamp 1620699047
<< nwell >>
rect -7185 2865 -7125 3110
<< poly >>
rect -5690 3235 -5650 3245
rect -5690 3215 -5680 3235
rect -5660 3215 -5650 3235
rect -5690 3205 -5650 3215
rect -7300 3130 -7120 3145
rect -7585 2850 -7545 2860
rect -7585 2830 -7575 2850
rect -7555 2830 -7545 2850
rect -7585 2820 -7545 2830
rect -7585 2435 -7570 2820
rect -5690 2555 -5675 3205
rect -3130 3190 -3010 3200
rect -3130 3170 -3120 3190
rect -3100 3185 -3010 3190
rect -3100 3170 -3090 3185
rect -3130 3160 -3090 3170
rect -7300 2540 -7120 2555
rect -6915 2540 -5675 2555
rect -7870 1730 -7830 1740
rect -7870 1710 -7860 1730
rect -7840 1710 -7830 1730
rect -7870 1700 -7830 1710
rect -3120 445 -3090 3160
rect -3060 2490 -3020 2500
rect -3060 2470 -3050 2490
rect -3030 2470 -3020 2490
rect -3060 2460 -3020 2470
rect 225 710 245 945
rect 225 700 265 710
rect 225 680 235 700
rect 255 680 265 700
rect 225 670 265 680
rect -3140 430 -3090 445
rect -3140 410 -3125 430
rect -3105 410 -3090 430
rect -3140 395 -3090 410
<< polycont >>
rect -5680 3215 -5660 3235
rect -7575 2830 -7555 2850
rect -3120 3170 -3100 3190
rect -7860 1710 -7840 1730
rect -3050 2470 -3030 2490
rect 235 680 255 700
rect -3125 410 -3105 430
<< locali >>
rect -5690 3260 -1300 3280
rect -5690 3235 -5650 3260
rect -5690 3215 -5680 3235
rect -5660 3215 -5650 3235
rect -5690 3205 -5650 3215
rect -1320 3210 -1300 3260
rect -3130 3190 -3090 3200
rect -1320 3190 0 3210
rect -3130 3185 -3120 3190
rect -7190 3170 -3120 3185
rect -3100 3170 -3090 3190
rect -7190 3165 -3090 3170
rect -7190 2860 -7165 3165
rect -3130 3160 -3090 3165
rect -5415 3020 -3040 3040
rect -7585 2850 -7510 2860
rect -7190 2855 -7115 2860
rect -7585 2830 -7575 2850
rect -7555 2830 -7510 2850
rect -7585 2820 -7510 2830
rect -7180 2820 -7115 2855
rect -6795 2820 -6770 2860
rect -6790 2520 -6770 2820
rect -5415 2560 -5395 3020
rect -5635 2540 -5395 2560
rect -5635 2520 -5615 2540
rect -7850 2500 -5615 2520
rect -3060 2500 -3040 3020
rect -7850 1740 -7830 2500
rect -3060 2490 -3020 2500
rect -3060 2470 -3050 2490
rect -3030 2470 -3020 2490
rect -3060 2460 -3020 2470
rect -7870 1730 -7830 1740
rect -7870 1710 -7860 1730
rect -7840 1710 -7830 1730
rect -7870 1700 -7830 1710
rect 135 765 185 1050
rect -155 730 8390 765
rect 225 700 265 710
rect 225 680 235 700
rect 255 680 265 700
rect 225 670 265 680
rect -3140 430 -3090 445
rect -3140 420 -3125 430
rect -4875 410 -3125 420
rect -3105 410 -3090 430
rect -4875 395 -3090 410
rect 8365 80 8390 730
rect 8365 75 8575 80
rect 8365 60 8580 75
<< viali >>
rect -7275 2905 -7245 2925
rect -6890 2905 -6860 2925
rect -7275 2750 -7245 2770
rect -6890 2750 -6860 2770
<< metal1 >>
rect -7290 2935 -6085 2940
rect -7290 2925 -6140 2935
rect -7290 2905 -7275 2925
rect -7245 2905 -6890 2925
rect -6860 2905 -6140 2925
rect -7290 2890 -6140 2905
rect -6145 2855 -6140 2890
rect -6090 2855 -6085 2935
rect -6145 2850 -6085 2855
rect -7290 2770 -6845 2785
rect -7290 2750 -7275 2770
rect -7245 2750 -6890 2770
rect -6860 2750 -6845 2770
rect -7290 2735 -6845 2750
rect -7165 2600 -7055 2735
rect -685 2660 10 2850
rect -7165 2330 -7060 2600
rect -190 2255 15 2445
rect -660 840 -465 925
rect 65 840 300 1180
rect -660 650 300 840
rect -5000 635 -4430 640
rect -5000 455 -4540 635
rect -4435 455 -4430 635
rect -5000 450 -4430 455
rect -660 365 -340 650
rect -5000 170 -340 365
<< via1 >>
rect -6140 2855 -6090 2935
rect -4540 455 -4435 635
<< metal2 >>
rect -6145 2935 -6085 2940
rect -6145 2855 -6140 2935
rect -6090 2855 -6085 2935
rect -6145 2330 -6085 2855
rect -2960 640 -2525 875
rect -1165 640 -730 875
rect -370 640 -190 1515
rect -4545 635 -190 640
rect -4545 455 -4540 635
rect -4435 615 -190 635
rect -4435 455 -200 615
rect -4545 450 -200 455
use adc_digital  adc_digital_0
timestamp 1620697130
transform 1 0 0 0 1 1665
box 0 -1665 25410 1645
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620697130
transform 1 0 -7585 0 1 -2490
box -255 2315 4445 5470
use comparator  comparator_0
timestamp 1620697130
transform 1 0 -2775 0 1 -1730
box -255 2315 2625 4970
use switch  switch_0
timestamp 1620697026
transform 1 0 -7425 0 1 2520
box -110 20 245 625
use switch  switch_1
timestamp 1620697026
transform 1 0 -7040 0 1 2520
box -110 20 245 625
<< end >>
