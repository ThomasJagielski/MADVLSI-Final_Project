magic
tech sky130A
timestamp 1620349204
<< end >>
