magic
tech sky130A
timestamp 1620670333
<< nwell >>
rect -120 155 410 395
<< nmos >>
rect 0 0 15 100
rect 65 0 80 100
rect 130 0 145 100
rect 195 0 210 100
rect 260 0 275 100
rect 325 0 340 100
<< pmos >>
rect 0 175 15 375
rect 65 175 80 375
rect 130 175 145 375
rect 195 175 210 375
rect 260 175 275 375
rect 325 175 340 375
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 145 85 195 100
rect 145 15 160 85
rect 180 15 195 85
rect 145 0 195 15
rect 210 85 260 100
rect 210 15 225 85
rect 245 15 260 85
rect 210 0 260 15
rect 275 85 325 100
rect 275 15 290 85
rect 310 15 325 85
rect 275 0 325 15
rect 340 85 390 100
rect 340 15 355 85
rect 375 15 390 85
rect 340 0 390 15
<< pdiff >>
rect -50 360 0 375
rect -50 190 -35 360
rect -15 190 0 360
rect -50 175 0 190
rect 15 360 65 375
rect 15 190 30 360
rect 50 190 65 360
rect 15 175 65 190
rect 80 360 130 375
rect 80 190 95 360
rect 115 190 130 360
rect 80 175 130 190
rect 145 360 195 375
rect 145 190 160 360
rect 180 190 195 360
rect 145 175 195 190
rect 210 360 260 375
rect 210 190 225 360
rect 245 190 260 360
rect 210 175 260 190
rect 275 360 325 375
rect 275 190 290 360
rect 310 190 325 360
rect 275 175 325 190
rect 340 360 390 375
rect 340 190 355 360
rect 375 190 390 360
rect 340 175 390 190
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
rect 160 15 180 85
rect 225 15 245 85
rect 290 15 310 85
rect 355 15 375 85
<< pdiffc >>
rect -35 190 -15 360
rect 30 190 50 360
rect 95 190 115 360
rect 160 190 180 360
rect 225 190 245 360
rect 290 190 310 360
rect 355 190 375 360
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 360 -50 375
rect -100 190 -85 360
rect -65 190 -50 360
rect -100 175 -50 190
<< psubdiffcont >>
rect -85 15 -65 85
<< nsubdiffcont >>
rect -85 190 -65 360
<< poly >>
rect 0 375 15 390
rect 65 375 80 390
rect 130 375 145 390
rect 195 375 210 390
rect 260 375 275 390
rect 325 375 340 390
rect 0 165 15 175
rect 65 165 80 175
rect 130 165 145 175
rect 195 165 210 175
rect 260 165 275 175
rect 325 165 340 175
rect 0 155 340 165
rect -70 150 340 155
rect -70 145 15 150
rect -70 125 -60 145
rect -40 125 15 145
rect -70 115 340 125
rect 0 110 340 115
rect 0 100 15 110
rect 65 100 80 110
rect 130 100 145 110
rect 195 100 210 110
rect 260 100 275 110
rect 325 100 340 110
rect 0 -15 15 0
rect 65 -15 80 0
rect 130 -15 145 0
rect 195 -15 210 0
rect 260 -15 275 0
rect 325 -15 340 0
<< polycont >>
rect -60 125 -40 145
<< locali >>
rect -50 390 385 410
rect -50 370 -5 390
rect -95 360 -5 370
rect -95 190 -85 360
rect -65 190 -35 360
rect -15 190 -5 360
rect -95 180 -5 190
rect 20 360 60 370
rect 20 190 30 360
rect 50 190 60 360
rect 20 160 60 190
rect 85 360 125 390
rect 85 190 95 360
rect 115 190 125 360
rect 85 180 125 190
rect 150 360 190 370
rect 150 190 160 360
rect 180 190 190 360
rect 150 160 190 190
rect 215 360 255 390
rect 215 190 225 360
rect 245 190 255 360
rect 215 180 255 190
rect 280 360 320 370
rect 280 190 290 360
rect 310 190 320 360
rect 280 160 320 190
rect 345 360 385 390
rect 345 190 355 360
rect 375 190 385 360
rect 345 180 385 190
rect -70 145 -30 155
rect -120 125 -60 145
rect -40 125 -30 145
rect -70 115 -30 125
rect 20 150 320 160
rect 20 125 410 150
rect 20 115 320 125
rect -95 85 -5 95
rect -95 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect -95 5 -5 15
rect 20 85 60 115
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect -45 -15 -5 5
rect 85 -15 125 15
rect 150 85 190 115
rect 150 15 160 85
rect 180 15 190 85
rect 150 5 190 15
rect 215 85 255 95
rect 215 15 225 85
rect 245 15 255 85
rect 215 -15 255 15
rect 280 85 320 115
rect 280 15 290 85
rect 310 15 320 85
rect 280 5 320 15
rect 345 85 385 95
rect 345 15 355 85
rect 375 15 385 85
rect 345 -15 385 15
rect -45 -35 385 -15
<< viali >>
rect -85 190 -65 360
rect -35 190 -15 360
rect 95 190 115 360
rect 225 190 245 360
rect 355 190 375 360
rect -85 15 -65 85
rect -35 15 -15 85
rect 95 15 115 85
rect 225 15 245 85
rect 355 15 375 85
<< metal1 >>
rect -120 360 410 370
rect -120 190 -85 360
rect -65 190 -35 360
rect -15 190 95 360
rect 115 190 225 360
rect 245 190 355 360
rect 375 190 410 360
rect -120 180 410 190
rect -120 85 410 95
rect -120 15 -85 85
rect -65 15 -35 85
rect -15 15 95 85
rect 115 15 225 85
rect 245 15 355 85
rect 375 15 410 85
rect -120 -100 410 15
<< labels >>
rlabel metal1 -120 275 -120 275 7 VDD
port 1 w
rlabel metal1 -120 -15 -120 -15 7 GND
port 2 w
rlabel locali -120 135 -120 135 7 A
port 3 w
rlabel locali 410 140 410 140 3 Y
port 4 e
<< end >>
