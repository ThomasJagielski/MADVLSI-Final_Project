magic
tech sky130A
timestamp 1620580153
<< nwell >>
rect -205 4650 2065 4900
rect 330 4530 435 4650
rect 1440 4620 1615 4650
rect 1440 4530 1545 4620
rect -205 3875 2065 4075
rect 340 3765 445 3875
rect 1420 3755 1525 3875
rect -205 2940 2065 3140
rect 215 2745 375 2940
rect 1360 2895 1855 2940
rect 1495 2745 1655 2895
<< nmos >>
rect -120 4345 -60 4495
rect 0 4345 60 4495
rect 120 4345 180 4495
rect 240 4345 300 4495
rect 360 4345 420 4495
rect 480 4345 540 4495
rect 600 4345 660 4495
rect 720 4345 780 4495
rect 840 4345 900 4495
rect 960 4345 1020 4495
rect 1080 4345 1140 4495
rect 1200 4345 1260 4495
rect 1320 4345 1380 4495
rect 1440 4345 1500 4495
rect 1560 4345 1620 4495
rect 1680 4345 1740 4495
rect 1800 4345 1860 4495
rect 1920 4345 1980 4495
rect -120 3460 -60 3610
rect 0 3460 60 3610
rect 120 3460 180 3610
rect 240 3460 300 3610
rect 360 3460 420 3610
rect 480 3460 540 3610
rect 600 3460 660 3610
rect 720 3460 780 3610
rect 840 3460 900 3610
rect 960 3460 1020 3610
rect 1080 3460 1140 3610
rect 1200 3460 1260 3610
rect 1320 3460 1380 3610
rect 1440 3460 1500 3610
rect 1560 3460 1620 3610
rect 1680 3460 1740 3610
rect 1800 3460 1860 3610
rect 1920 3460 1980 3610
rect -120 2430 -60 2580
rect 0 2430 60 2580
rect 120 2430 180 2580
rect 240 2430 300 2580
rect 360 2430 420 2580
rect 480 2430 540 2580
rect 600 2430 660 2580
rect 720 2430 780 2580
rect 840 2430 900 2580
rect 960 2430 1020 2580
rect 1080 2430 1140 2580
rect 1200 2430 1260 2580
rect 1320 2430 1380 2580
rect 1440 2430 1500 2580
rect 1560 2430 1620 2580
rect 1680 2430 1740 2580
rect 1800 2430 1860 2580
rect 1920 2430 1980 2580
<< pmos >>
rect -120 4675 -60 4825
rect 0 4675 60 4825
rect 120 4675 180 4825
rect 240 4675 300 4825
rect 360 4675 420 4825
rect 480 4675 540 4825
rect 600 4675 660 4825
rect 720 4675 780 4825
rect 840 4675 900 4825
rect 960 4675 1020 4825
rect 1080 4675 1140 4825
rect 1200 4675 1260 4825
rect 1320 4675 1380 4825
rect 1440 4675 1500 4825
rect 1560 4675 1620 4825
rect 1680 4675 1740 4825
rect 1800 4675 1860 4825
rect 1920 4675 1980 4825
rect -120 3900 -60 4050
rect 0 3900 60 4050
rect 120 3900 180 4050
rect 240 3900 300 4050
rect 360 3900 420 4050
rect 480 3900 540 4050
rect 600 3900 660 4050
rect 720 3900 780 4050
rect 840 3900 900 4050
rect 960 3900 1020 4050
rect 1080 3900 1140 4050
rect 1200 3900 1260 4050
rect 1320 3900 1380 4050
rect 1440 3900 1500 4050
rect 1560 3900 1620 4050
rect 1680 3900 1740 4050
rect 1800 3900 1860 4050
rect 1920 3900 1980 4050
rect -120 2965 -60 3115
rect 0 2965 60 3115
rect 120 2965 180 3115
rect 240 2965 300 3115
rect 360 2965 420 3115
rect 480 2965 540 3115
rect 600 2965 660 3115
rect 720 2965 780 3115
rect 840 2965 900 3115
rect 960 2965 1020 3115
rect 1080 2965 1140 3115
rect 1200 2965 1260 3115
rect 1320 2965 1380 3115
rect 1440 2965 1500 3115
rect 1560 2965 1620 3115
rect 1680 2965 1740 3115
rect 1800 2965 1860 3115
rect 1920 2965 1980 3115
<< ndiff >>
rect -180 4480 -120 4495
rect -180 4360 -165 4480
rect -135 4360 -120 4480
rect -180 4345 -120 4360
rect -60 4480 0 4495
rect -60 4360 -45 4480
rect -15 4360 0 4480
rect -60 4345 0 4360
rect 60 4480 120 4495
rect 60 4360 75 4480
rect 105 4360 120 4480
rect 60 4345 120 4360
rect 180 4480 240 4495
rect 180 4360 195 4480
rect 225 4360 240 4480
rect 180 4345 240 4360
rect 300 4480 360 4495
rect 300 4360 315 4480
rect 345 4360 360 4480
rect 300 4345 360 4360
rect 420 4480 480 4495
rect 420 4360 435 4480
rect 465 4360 480 4480
rect 420 4345 480 4360
rect 540 4480 600 4495
rect 540 4360 555 4480
rect 585 4360 600 4480
rect 540 4345 600 4360
rect 660 4480 720 4495
rect 660 4360 675 4480
rect 705 4360 720 4480
rect 660 4345 720 4360
rect 780 4480 840 4495
rect 780 4360 795 4480
rect 825 4360 840 4480
rect 780 4345 840 4360
rect 900 4480 960 4495
rect 900 4360 915 4480
rect 945 4360 960 4480
rect 900 4345 960 4360
rect 1020 4480 1080 4495
rect 1020 4360 1035 4480
rect 1065 4360 1080 4480
rect 1020 4345 1080 4360
rect 1140 4480 1200 4495
rect 1140 4360 1155 4480
rect 1185 4360 1200 4480
rect 1140 4345 1200 4360
rect 1260 4480 1320 4495
rect 1260 4360 1275 4480
rect 1305 4360 1320 4480
rect 1260 4345 1320 4360
rect 1380 4480 1440 4495
rect 1380 4360 1395 4480
rect 1425 4360 1440 4480
rect 1380 4345 1440 4360
rect 1500 4480 1560 4495
rect 1500 4360 1515 4480
rect 1545 4360 1560 4480
rect 1500 4345 1560 4360
rect 1620 4480 1680 4495
rect 1620 4360 1635 4480
rect 1665 4360 1680 4480
rect 1620 4345 1680 4360
rect 1740 4480 1800 4495
rect 1740 4360 1755 4480
rect 1785 4360 1800 4480
rect 1740 4345 1800 4360
rect 1860 4480 1920 4495
rect 1860 4360 1875 4480
rect 1905 4360 1920 4480
rect 1860 4345 1920 4360
rect 1980 4480 2040 4495
rect 1980 4360 1995 4480
rect 2025 4360 2040 4480
rect 1980 4345 2040 4360
rect -180 3595 -120 3610
rect -180 3475 -165 3595
rect -135 3475 -120 3595
rect -180 3460 -120 3475
rect -60 3595 0 3610
rect -60 3475 -45 3595
rect -15 3475 0 3595
rect -60 3460 0 3475
rect 60 3595 120 3610
rect 60 3475 75 3595
rect 105 3475 120 3595
rect 60 3460 120 3475
rect 180 3595 240 3610
rect 180 3475 195 3595
rect 225 3475 240 3595
rect 180 3460 240 3475
rect 300 3595 360 3610
rect 300 3475 315 3595
rect 345 3475 360 3595
rect 300 3460 360 3475
rect 420 3595 480 3610
rect 420 3475 435 3595
rect 465 3475 480 3595
rect 420 3460 480 3475
rect 540 3595 600 3610
rect 540 3475 555 3595
rect 585 3475 600 3595
rect 540 3460 600 3475
rect 660 3595 720 3610
rect 660 3475 675 3595
rect 705 3475 720 3595
rect 660 3460 720 3475
rect 780 3595 840 3610
rect 780 3475 795 3595
rect 825 3475 840 3595
rect 780 3460 840 3475
rect 900 3595 960 3610
rect 900 3475 915 3595
rect 945 3475 960 3595
rect 900 3460 960 3475
rect 1020 3595 1080 3610
rect 1020 3475 1035 3595
rect 1065 3475 1080 3595
rect 1020 3460 1080 3475
rect 1140 3595 1200 3610
rect 1140 3475 1155 3595
rect 1185 3475 1200 3595
rect 1140 3460 1200 3475
rect 1260 3595 1320 3610
rect 1260 3475 1275 3595
rect 1305 3475 1320 3595
rect 1260 3460 1320 3475
rect 1380 3595 1440 3610
rect 1380 3475 1395 3595
rect 1425 3475 1440 3595
rect 1380 3460 1440 3475
rect 1500 3595 1560 3610
rect 1500 3475 1515 3595
rect 1545 3475 1560 3595
rect 1500 3460 1560 3475
rect 1620 3595 1680 3610
rect 1620 3475 1635 3595
rect 1665 3475 1680 3595
rect 1620 3460 1680 3475
rect 1740 3595 1800 3610
rect 1740 3475 1755 3595
rect 1785 3475 1800 3595
rect 1740 3460 1800 3475
rect 1860 3595 1920 3610
rect 1860 3475 1875 3595
rect 1905 3475 1920 3595
rect 1860 3460 1920 3475
rect 1980 3595 2040 3610
rect 1980 3475 1995 3595
rect 2025 3475 2040 3595
rect 1980 3460 2040 3475
rect -180 2565 -120 2580
rect -180 2445 -165 2565
rect -135 2445 -120 2565
rect -180 2430 -120 2445
rect -60 2565 0 2580
rect -60 2445 -45 2565
rect -15 2445 0 2565
rect -60 2430 0 2445
rect 60 2565 120 2580
rect 60 2445 75 2565
rect 105 2445 120 2565
rect 60 2430 120 2445
rect 180 2565 240 2580
rect 180 2445 195 2565
rect 225 2445 240 2565
rect 180 2430 240 2445
rect 300 2565 360 2580
rect 300 2445 315 2565
rect 345 2445 360 2565
rect 300 2430 360 2445
rect 420 2565 480 2580
rect 420 2445 435 2565
rect 465 2445 480 2565
rect 420 2430 480 2445
rect 540 2565 600 2580
rect 540 2445 555 2565
rect 585 2445 600 2565
rect 540 2430 600 2445
rect 660 2565 720 2580
rect 660 2445 675 2565
rect 705 2445 720 2565
rect 660 2430 720 2445
rect 780 2565 840 2580
rect 780 2445 795 2565
rect 825 2445 840 2565
rect 780 2430 840 2445
rect 900 2565 960 2580
rect 900 2445 915 2565
rect 945 2445 960 2565
rect 900 2430 960 2445
rect 1020 2565 1080 2580
rect 1020 2445 1035 2565
rect 1065 2445 1080 2565
rect 1020 2430 1080 2445
rect 1140 2565 1200 2580
rect 1140 2445 1155 2565
rect 1185 2445 1200 2565
rect 1140 2430 1200 2445
rect 1260 2565 1320 2580
rect 1260 2445 1275 2565
rect 1305 2445 1320 2565
rect 1260 2430 1320 2445
rect 1380 2565 1440 2580
rect 1380 2445 1395 2565
rect 1425 2445 1440 2565
rect 1380 2430 1440 2445
rect 1500 2565 1560 2580
rect 1500 2445 1515 2565
rect 1545 2445 1560 2565
rect 1500 2430 1560 2445
rect 1620 2565 1680 2580
rect 1620 2445 1635 2565
rect 1665 2445 1680 2565
rect 1620 2430 1680 2445
rect 1740 2565 1800 2580
rect 1740 2445 1755 2565
rect 1785 2445 1800 2565
rect 1740 2430 1800 2445
rect 1860 2565 1920 2580
rect 1860 2445 1875 2565
rect 1905 2445 1920 2565
rect 1860 2430 1920 2445
rect 1980 2565 2040 2580
rect 1980 2445 1995 2565
rect 2025 2445 2040 2565
rect 1980 2430 2040 2445
<< pdiff >>
rect -180 4810 -120 4825
rect -180 4690 -165 4810
rect -135 4690 -120 4810
rect -180 4675 -120 4690
rect -60 4810 0 4825
rect -60 4690 -45 4810
rect -15 4690 0 4810
rect -60 4675 0 4690
rect 60 4810 120 4825
rect 60 4690 75 4810
rect 105 4690 120 4810
rect 60 4675 120 4690
rect 180 4810 240 4825
rect 180 4690 195 4810
rect 225 4690 240 4810
rect 180 4675 240 4690
rect 300 4810 360 4825
rect 300 4690 315 4810
rect 345 4690 360 4810
rect 300 4675 360 4690
rect 420 4810 480 4825
rect 420 4690 435 4810
rect 465 4690 480 4810
rect 420 4675 480 4690
rect 540 4810 600 4825
rect 540 4690 555 4810
rect 585 4690 600 4810
rect 540 4675 600 4690
rect 660 4810 720 4825
rect 660 4690 675 4810
rect 705 4690 720 4810
rect 660 4675 720 4690
rect 780 4810 840 4825
rect 780 4690 795 4810
rect 825 4690 840 4810
rect 780 4675 840 4690
rect 900 4810 960 4825
rect 900 4690 915 4810
rect 945 4690 960 4810
rect 900 4675 960 4690
rect 1020 4810 1080 4825
rect 1020 4690 1035 4810
rect 1065 4690 1080 4810
rect 1020 4675 1080 4690
rect 1140 4810 1200 4825
rect 1140 4690 1155 4810
rect 1185 4690 1200 4810
rect 1140 4675 1200 4690
rect 1260 4810 1320 4825
rect 1260 4690 1275 4810
rect 1305 4690 1320 4810
rect 1260 4675 1320 4690
rect 1380 4810 1440 4825
rect 1380 4690 1395 4810
rect 1425 4690 1440 4810
rect 1380 4675 1440 4690
rect 1500 4810 1560 4825
rect 1500 4690 1515 4810
rect 1545 4690 1560 4810
rect 1500 4675 1560 4690
rect 1620 4810 1680 4825
rect 1620 4690 1635 4810
rect 1665 4690 1680 4810
rect 1620 4675 1680 4690
rect 1740 4810 1800 4825
rect 1740 4690 1755 4810
rect 1785 4690 1800 4810
rect 1740 4675 1800 4690
rect 1860 4810 1920 4825
rect 1860 4690 1875 4810
rect 1905 4690 1920 4810
rect 1860 4675 1920 4690
rect 1980 4810 2040 4825
rect 1980 4690 1995 4810
rect 2025 4690 2040 4810
rect 1980 4675 2040 4690
rect -180 4035 -120 4050
rect -180 3915 -165 4035
rect -135 3915 -120 4035
rect -180 3900 -120 3915
rect -60 4035 0 4050
rect -60 3915 -45 4035
rect -15 3915 0 4035
rect -60 3900 0 3915
rect 60 4035 120 4050
rect 60 3915 75 4035
rect 105 3915 120 4035
rect 60 3900 120 3915
rect 180 4035 240 4050
rect 180 3915 195 4035
rect 225 3915 240 4035
rect 180 3900 240 3915
rect 300 4035 360 4050
rect 300 3915 315 4035
rect 345 3915 360 4035
rect 300 3900 360 3915
rect 420 4035 480 4050
rect 420 3915 435 4035
rect 465 3915 480 4035
rect 420 3900 480 3915
rect 540 4035 600 4050
rect 540 3915 555 4035
rect 585 3915 600 4035
rect 540 3900 600 3915
rect 660 4035 720 4050
rect 660 3915 675 4035
rect 705 3915 720 4035
rect 660 3900 720 3915
rect 780 4035 840 4050
rect 780 3915 795 4035
rect 825 3915 840 4035
rect 780 3900 840 3915
rect 900 4035 960 4050
rect 900 3915 915 4035
rect 945 3915 960 4035
rect 900 3900 960 3915
rect 1020 4035 1080 4050
rect 1020 3915 1035 4035
rect 1065 3915 1080 4035
rect 1020 3900 1080 3915
rect 1140 4035 1200 4050
rect 1140 3915 1155 4035
rect 1185 3915 1200 4035
rect 1140 3900 1200 3915
rect 1260 4035 1320 4050
rect 1260 3915 1275 4035
rect 1305 3915 1320 4035
rect 1260 3900 1320 3915
rect 1380 4035 1440 4050
rect 1380 3915 1395 4035
rect 1425 3915 1440 4035
rect 1380 3900 1440 3915
rect 1500 4035 1560 4050
rect 1500 3915 1515 4035
rect 1545 3915 1560 4035
rect 1500 3900 1560 3915
rect 1620 4035 1680 4050
rect 1620 3915 1635 4035
rect 1665 3915 1680 4035
rect 1620 3900 1680 3915
rect 1740 4035 1800 4050
rect 1740 3915 1755 4035
rect 1785 3915 1800 4035
rect 1740 3900 1800 3915
rect 1860 4035 1920 4050
rect 1860 3915 1875 4035
rect 1905 3915 1920 4035
rect 1860 3900 1920 3915
rect 1980 4035 2040 4050
rect 1980 3915 1995 4035
rect 2025 3915 2040 4035
rect 1980 3900 2040 3915
rect -180 3100 -120 3115
rect -180 2980 -165 3100
rect -135 2980 -120 3100
rect -180 2965 -120 2980
rect -60 3100 0 3115
rect -60 2980 -45 3100
rect -15 2980 0 3100
rect -60 2965 0 2980
rect 60 3100 120 3115
rect 60 2980 75 3100
rect 105 2980 120 3100
rect 60 2965 120 2980
rect 180 3100 240 3115
rect 180 2980 195 3100
rect 225 2980 240 3100
rect 180 2965 240 2980
rect 300 3100 360 3115
rect 300 2980 315 3100
rect 345 2980 360 3100
rect 300 2965 360 2980
rect 420 3100 480 3115
rect 420 2980 435 3100
rect 465 2980 480 3100
rect 420 2965 480 2980
rect 540 3100 600 3115
rect 540 2980 555 3100
rect 585 2980 600 3100
rect 540 2965 600 2980
rect 660 3100 720 3115
rect 660 2980 675 3100
rect 705 2980 720 3100
rect 660 2965 720 2980
rect 780 3100 840 3115
rect 780 2980 795 3100
rect 825 2980 840 3100
rect 780 2965 840 2980
rect 900 3100 960 3115
rect 900 2980 915 3100
rect 945 2980 960 3100
rect 900 2965 960 2980
rect 1020 3100 1080 3115
rect 1020 2980 1035 3100
rect 1065 2980 1080 3100
rect 1020 2965 1080 2980
rect 1140 3100 1200 3115
rect 1140 2980 1155 3100
rect 1185 2980 1200 3100
rect 1140 2965 1200 2980
rect 1260 3100 1320 3115
rect 1260 2980 1275 3100
rect 1305 2980 1320 3100
rect 1260 2965 1320 2980
rect 1380 3100 1440 3115
rect 1380 2980 1395 3100
rect 1425 2980 1440 3100
rect 1380 2965 1440 2980
rect 1500 3100 1560 3115
rect 1500 2980 1515 3100
rect 1545 2980 1560 3100
rect 1500 2965 1560 2980
rect 1620 3100 1680 3115
rect 1620 2980 1635 3100
rect 1665 2980 1680 3100
rect 1620 2965 1680 2980
rect 1740 3100 1800 3115
rect 1740 2980 1755 3100
rect 1785 2980 1800 3100
rect 1740 2965 1800 2980
rect 1860 3100 1920 3115
rect 1860 2980 1875 3100
rect 1905 2980 1920 3100
rect 1860 2965 1920 2980
rect 1980 3100 2040 3115
rect 1980 2980 1995 3100
rect 2025 2980 2040 3100
rect 1980 2965 2040 2980
<< ndiffc >>
rect -165 4360 -135 4480
rect -45 4360 -15 4480
rect 75 4360 105 4480
rect 195 4360 225 4480
rect 315 4360 345 4480
rect 435 4360 465 4480
rect 555 4360 585 4480
rect 675 4360 705 4480
rect 795 4360 825 4480
rect 915 4360 945 4480
rect 1035 4360 1065 4480
rect 1155 4360 1185 4480
rect 1275 4360 1305 4480
rect 1395 4360 1425 4480
rect 1515 4360 1545 4480
rect 1635 4360 1665 4480
rect 1755 4360 1785 4480
rect 1875 4360 1905 4480
rect 1995 4360 2025 4480
rect -165 3475 -135 3595
rect -45 3475 -15 3595
rect 75 3475 105 3595
rect 195 3475 225 3595
rect 315 3475 345 3595
rect 435 3475 465 3595
rect 555 3475 585 3595
rect 675 3475 705 3595
rect 795 3475 825 3595
rect 915 3475 945 3595
rect 1035 3475 1065 3595
rect 1155 3475 1185 3595
rect 1275 3475 1305 3595
rect 1395 3475 1425 3595
rect 1515 3475 1545 3595
rect 1635 3475 1665 3595
rect 1755 3475 1785 3595
rect 1875 3475 1905 3595
rect 1995 3475 2025 3595
rect -165 2445 -135 2565
rect -45 2445 -15 2565
rect 75 2445 105 2565
rect 195 2445 225 2565
rect 315 2445 345 2565
rect 435 2445 465 2565
rect 555 2445 585 2565
rect 675 2445 705 2565
rect 795 2445 825 2565
rect 915 2445 945 2565
rect 1035 2445 1065 2565
rect 1155 2445 1185 2565
rect 1275 2445 1305 2565
rect 1395 2445 1425 2565
rect 1515 2445 1545 2565
rect 1635 2445 1665 2565
rect 1755 2445 1785 2565
rect 1875 2445 1905 2565
rect 1995 2445 2025 2565
<< pdiffc >>
rect -165 4690 -135 4810
rect -45 4690 -15 4810
rect 75 4690 105 4810
rect 195 4690 225 4810
rect 315 4690 345 4810
rect 435 4690 465 4810
rect 555 4690 585 4810
rect 675 4690 705 4810
rect 795 4690 825 4810
rect 915 4690 945 4810
rect 1035 4690 1065 4810
rect 1155 4690 1185 4810
rect 1275 4690 1305 4810
rect 1395 4690 1425 4810
rect 1515 4690 1545 4810
rect 1635 4690 1665 4810
rect 1755 4690 1785 4810
rect 1875 4690 1905 4810
rect 1995 4690 2025 4810
rect -165 3915 -135 4035
rect -45 3915 -15 4035
rect 75 3915 105 4035
rect 195 3915 225 4035
rect 315 3915 345 4035
rect 435 3915 465 4035
rect 555 3915 585 4035
rect 675 3915 705 4035
rect 795 3915 825 4035
rect 915 3915 945 4035
rect 1035 3915 1065 4035
rect 1155 3915 1185 4035
rect 1275 3915 1305 4035
rect 1395 3915 1425 4035
rect 1515 3915 1545 4035
rect 1635 3915 1665 4035
rect 1755 3915 1785 4035
rect 1875 3915 1905 4035
rect 1995 3915 2025 4035
rect -165 2980 -135 3100
rect -45 2980 -15 3100
rect 75 2980 105 3100
rect 195 2980 225 3100
rect 315 2980 345 3100
rect 435 2980 465 3100
rect 555 2980 585 3100
rect 675 2980 705 3100
rect 795 2980 825 3100
rect 915 2980 945 3100
rect 1035 2980 1065 3100
rect 1155 2980 1185 3100
rect 1275 2980 1305 3100
rect 1395 2980 1425 3100
rect 1515 2980 1545 3100
rect 1635 2980 1665 3100
rect 1755 2980 1785 3100
rect 1875 2980 1905 3100
rect 1995 2980 2025 3100
<< psubdiff >>
rect 165 4575 225 4590
rect 165 4545 180 4575
rect 210 4545 225 4575
rect 165 4530 225 4545
rect 1720 4590 1780 4605
rect 1720 4560 1735 4590
rect 1765 4560 1780 4590
rect 1720 4545 1780 4560
rect 165 3755 225 3770
rect 165 3720 180 3755
rect 210 3720 225 3755
rect 1675 3745 1735 3760
rect 165 3705 225 3720
rect 1675 3710 1690 3745
rect 1720 3710 1735 3745
rect 1675 3695 1735 3710
rect 450 2730 570 2745
rect 450 2640 465 2730
rect 555 2640 570 2730
rect 1290 2730 1410 2745
rect 450 2625 570 2640
rect 1290 2640 1305 2730
rect 1395 2640 1410 2730
rect 1290 2625 1410 2640
<< nsubdiff >>
rect 350 4595 410 4605
rect 350 4565 365 4595
rect 395 4565 410 4595
rect 350 4550 410 4565
rect 1460 4595 1520 4605
rect 1460 4565 1475 4595
rect 1505 4565 1520 4595
rect 1460 4550 1520 4565
rect 360 3835 420 3850
rect 360 3800 375 3835
rect 405 3800 420 3835
rect 1440 3825 1500 3840
rect 360 3785 420 3800
rect 1440 3790 1455 3825
rect 1485 3790 1500 3825
rect 1440 3775 1500 3790
rect 235 2870 355 2885
rect 235 2780 250 2870
rect 340 2780 355 2870
rect 1515 2870 1635 2885
rect 235 2765 355 2780
rect 1515 2780 1530 2870
rect 1620 2780 1635 2870
rect 1515 2765 1635 2780
<< psubdiffcont >>
rect 180 4545 210 4575
rect 1735 4560 1765 4590
rect 180 3720 210 3755
rect 1690 3710 1720 3745
rect 465 2640 555 2730
rect 1305 2640 1395 2730
<< nsubdiffcont >>
rect 365 4565 395 4595
rect 1475 4565 1505 4595
rect 375 3800 405 3835
rect 1455 3790 1485 3825
rect 250 2780 340 2870
rect 1530 2780 1620 2870
<< poly >>
rect -240 4915 1380 4930
rect -120 4825 -60 4840
rect 0 4825 60 4840
rect 120 4825 180 4840
rect 240 4825 300 4840
rect 360 4825 420 4840
rect 480 4825 540 4915
rect 615 4870 655 4880
rect 615 4850 625 4870
rect 645 4850 655 4870
rect 615 4840 655 4850
rect 1200 4870 1240 4880
rect 1200 4850 1210 4870
rect 1230 4850 1240 4870
rect 1200 4840 1240 4850
rect 600 4825 660 4840
rect 720 4825 780 4840
rect 840 4825 900 4840
rect 960 4825 1020 4840
rect 1080 4825 1140 4840
rect 1200 4825 1260 4840
rect 1320 4825 1380 4915
rect 1440 4825 1500 4840
rect 1560 4825 1620 4840
rect 1680 4825 1740 4840
rect 1800 4825 1860 4840
rect 1920 4825 1980 4840
rect -120 4660 -60 4675
rect 0 4660 60 4675
rect 120 4660 180 4675
rect 240 4660 300 4675
rect 360 4660 420 4675
rect -175 4650 420 4660
rect -175 4630 -165 4650
rect -70 4630 -45 4650
rect 50 4630 75 4650
rect 170 4630 195 4650
rect 290 4630 315 4650
rect 410 4630 420 4650
rect -175 4620 420 4630
rect -120 4495 -60 4510
rect 0 4495 60 4510
rect 120 4495 180 4510
rect 240 4495 300 4510
rect 360 4495 420 4510
rect 480 4495 540 4675
rect 600 4660 660 4675
rect 720 4635 780 4675
rect 600 4620 780 4635
rect 600 4495 660 4620
rect 840 4590 900 4675
rect 960 4590 1020 4675
rect 1080 4635 1140 4675
rect 1200 4660 1260 4675
rect 1080 4620 1260 4635
rect 840 4580 1020 4590
rect 840 4575 920 4580
rect 910 4560 920 4575
rect 940 4575 1020 4580
rect 940 4560 950 4575
rect 910 4550 950 4560
rect 720 4495 780 4510
rect 840 4495 900 4510
rect 960 4495 1020 4510
rect 1080 4495 1140 4510
rect 1200 4495 1260 4620
rect 1320 4495 1380 4675
rect 1440 4660 1500 4675
rect 1560 4660 1620 4675
rect 1680 4660 1740 4675
rect 1800 4660 1860 4675
rect 1920 4660 1980 4675
rect 1440 4650 2035 4660
rect 1440 4630 1450 4650
rect 1545 4630 1570 4650
rect 1665 4630 1690 4650
rect 1785 4630 1810 4650
rect 1905 4630 1930 4650
rect 2025 4630 2035 4650
rect 1440 4620 2035 4630
rect 2020 4540 2060 4550
rect 2020 4520 2030 4540
rect 2050 4525 2060 4540
rect 2050 4520 2075 4525
rect 2020 4510 2075 4520
rect 1440 4495 1500 4510
rect 1560 4495 1620 4510
rect 1680 4495 1740 4510
rect 1800 4495 1860 4510
rect 1920 4495 1980 4510
rect -120 4330 -60 4345
rect 0 4330 60 4345
rect 120 4330 180 4345
rect 240 4330 300 4345
rect 360 4330 420 4345
rect 480 4330 540 4345
rect -175 4320 420 4330
rect -175 4300 -165 4320
rect -70 4300 -45 4320
rect 50 4300 75 4320
rect 170 4300 195 4320
rect 290 4300 315 4320
rect 410 4300 420 4320
rect -175 4290 420 4300
rect 600 4205 660 4345
rect 720 4330 780 4345
rect 725 4325 765 4330
rect 725 4305 735 4325
rect 755 4305 765 4325
rect 725 4295 765 4305
rect 840 4305 900 4345
rect 960 4305 1020 4345
rect 1080 4330 1140 4345
rect 1200 4330 1260 4345
rect 1320 4330 1380 4345
rect 1440 4330 1500 4345
rect 1560 4330 1620 4345
rect 1680 4330 1740 4345
rect 1800 4330 1860 4345
rect 1920 4330 1980 4345
rect -240 4190 660 4205
rect 840 4290 1020 4305
rect 1095 4325 1135 4330
rect 1095 4305 1105 4325
rect 1125 4305 1135 4325
rect 1095 4295 1135 4305
rect 1440 4320 2035 4330
rect 1440 4300 1450 4320
rect 1545 4300 1570 4320
rect 1665 4300 1690 4320
rect 1785 4300 1810 4320
rect 1905 4300 1930 4320
rect 2025 4300 2035 4320
rect 1440 4290 2035 4300
rect 840 4165 855 4290
rect -220 4150 855 4165
rect -220 3690 -205 4150
rect 2060 4105 2075 4510
rect 360 4090 2075 4105
rect -120 4050 -60 4065
rect 0 4050 60 4065
rect 120 4050 180 4065
rect 240 4050 300 4065
rect 360 4050 420 4090
rect 480 4050 540 4065
rect 600 4050 660 4065
rect 720 4050 780 4090
rect 840 4050 900 4065
rect 960 4050 1020 4065
rect 1080 4050 1140 4090
rect 1200 4050 1260 4065
rect 1320 4050 1380 4065
rect 1440 4050 1500 4090
rect 1560 4050 1620 4065
rect 1680 4050 1740 4065
rect 1800 4050 1860 4065
rect 1920 4050 1980 4065
rect -120 3885 -60 3900
rect 0 3885 60 3900
rect 120 3885 180 3900
rect 240 3885 300 3900
rect 360 3885 420 3900
rect -175 3875 300 3885
rect -175 3855 -165 3875
rect -70 3855 -45 3875
rect 50 3855 75 3875
rect 170 3855 195 3875
rect 290 3855 300 3875
rect -175 3845 300 3855
rect 480 3875 540 3900
rect 600 3885 660 3900
rect 720 3885 780 3900
rect 480 3855 490 3875
rect 530 3855 540 3875
rect 480 3845 540 3855
rect 620 3875 660 3885
rect 620 3855 630 3875
rect 650 3855 660 3875
rect 620 3845 660 3855
rect 840 3875 900 3900
rect 840 3855 850 3875
rect 890 3855 900 3875
rect 840 3845 900 3855
rect 960 3875 1020 3900
rect 1080 3885 1140 3900
rect 1200 3885 1260 3900
rect 960 3855 970 3875
rect 1010 3855 1020 3875
rect 960 3845 1020 3855
rect 1200 3875 1240 3885
rect 1200 3855 1210 3875
rect 1230 3855 1240 3875
rect 1200 3845 1240 3855
rect 1320 3875 1380 3900
rect 1440 3885 1500 3900
rect 1560 3885 1620 3900
rect 1680 3885 1740 3900
rect 1800 3885 1860 3900
rect 1920 3885 1980 3900
rect 1320 3855 1330 3875
rect 1370 3855 1380 3875
rect 1320 3845 1380 3855
rect 1560 3875 2035 3885
rect 1560 3855 1570 3875
rect 1665 3855 1690 3875
rect 1785 3855 1810 3875
rect 1905 3855 1930 3875
rect 2025 3855 2035 3875
rect 1560 3845 2035 3855
rect 910 3815 950 3825
rect 910 3795 920 3815
rect 940 3795 950 3815
rect 910 3785 950 3795
rect 920 3725 940 3785
rect 910 3715 950 3725
rect 910 3695 920 3715
rect 940 3695 950 3715
rect -220 3675 420 3690
rect 910 3685 950 3695
rect -120 3610 -60 3625
rect 0 3610 60 3625
rect 120 3610 180 3625
rect 240 3610 300 3625
rect 360 3610 420 3675
rect 480 3655 540 3665
rect 480 3635 490 3655
rect 530 3635 540 3655
rect 480 3610 540 3635
rect 620 3655 660 3665
rect 620 3635 630 3655
rect 650 3635 660 3655
rect 620 3625 660 3635
rect 840 3655 900 3665
rect 840 3635 850 3655
rect 890 3635 900 3655
rect 600 3610 660 3625
rect 720 3610 780 3625
rect 840 3610 900 3635
rect 960 3655 1020 3665
rect 960 3635 970 3655
rect 1010 3635 1020 3655
rect 960 3610 1020 3635
rect 1200 3655 1240 3665
rect 1200 3635 1210 3655
rect 1230 3635 1240 3655
rect 1200 3625 1240 3635
rect 1320 3655 1380 3665
rect 1320 3635 1330 3655
rect 1370 3635 1380 3655
rect 1080 3610 1140 3625
rect 1200 3610 1260 3625
rect 1320 3610 1380 3635
rect 1440 3610 1500 3625
rect 1560 3610 1620 3625
rect 1680 3610 1740 3625
rect 1800 3610 1860 3625
rect 1920 3610 1980 3625
rect -120 3445 -60 3460
rect 0 3445 60 3460
rect 120 3445 180 3460
rect 240 3445 300 3460
rect -175 3435 300 3445
rect -175 3415 -165 3435
rect -70 3415 -45 3435
rect 50 3415 75 3435
rect 170 3415 195 3435
rect 290 3415 300 3435
rect -175 3405 300 3415
rect 360 3420 420 3460
rect 480 3445 540 3460
rect 600 3445 660 3460
rect 720 3420 780 3460
rect 840 3445 900 3460
rect 960 3445 1020 3460
rect 1080 3420 1140 3460
rect 1200 3445 1260 3460
rect 1320 3445 1380 3460
rect 1440 3420 1500 3460
rect 360 3405 1500 3420
rect 1560 3445 1620 3460
rect 1680 3445 1740 3460
rect 1800 3445 1860 3460
rect 1920 3445 1980 3460
rect 1560 3435 2035 3445
rect 1560 3415 1570 3435
rect 1665 3415 1690 3435
rect 1785 3415 1810 3435
rect 1905 3415 1930 3435
rect 2025 3415 2035 3435
rect 1560 3405 2035 3415
rect 440 3190 460 3405
rect 360 3180 400 3190
rect 360 3160 370 3180
rect 390 3160 400 3180
rect 360 3130 400 3160
rect 430 3180 470 3190
rect 430 3160 440 3180
rect 460 3160 470 3180
rect 430 3150 470 3160
rect 720 3180 760 3190
rect 720 3160 730 3180
rect 750 3160 760 3180
rect 720 3130 760 3160
rect 1100 3180 1140 3190
rect 1100 3160 1110 3180
rect 1130 3160 1140 3180
rect 1100 3130 1140 3160
rect 1460 3180 1500 3190
rect 1460 3160 1470 3180
rect 1490 3160 1500 3180
rect 2060 3175 2075 4090
rect 1460 3130 1500 3160
rect 1800 3160 2075 3175
rect -120 3115 -60 3130
rect 0 3115 60 3130
rect 120 3115 180 3130
rect 240 3115 300 3130
rect 360 3115 420 3130
rect 480 3115 540 3130
rect 600 3115 660 3130
rect 720 3115 780 3130
rect 840 3115 900 3130
rect 960 3115 1020 3130
rect 1080 3115 1140 3130
rect 1200 3115 1260 3130
rect 1320 3115 1380 3130
rect 1440 3115 1500 3130
rect 1560 3115 1620 3130
rect 1680 3115 1740 3130
rect 1800 3115 1860 3160
rect 1920 3115 1980 3130
rect -120 2950 -60 2965
rect -175 2940 -60 2950
rect -175 2920 -165 2940
rect -70 2920 -60 2940
rect -175 2910 -60 2920
rect 0 2925 60 2965
rect 120 2925 180 2965
rect 240 2925 300 2965
rect 360 2950 420 2965
rect 480 2925 540 2965
rect 600 2925 660 2965
rect 720 2950 780 2965
rect 840 2925 900 2965
rect 960 2925 1020 2965
rect 1080 2950 1140 2965
rect 1200 2925 1260 2965
rect 1320 2925 1380 2965
rect 1440 2950 1500 2965
rect 1560 2925 1620 2965
rect 1680 2925 1740 2965
rect 1800 2925 1860 2965
rect 0 2910 1860 2925
rect 1920 2950 1980 2965
rect 1920 2940 2035 2950
rect 1920 2920 1930 2940
rect 2025 2920 2035 2940
rect 1920 2910 2035 2920
rect 785 2875 835 2885
rect 785 2850 795 2875
rect 825 2855 835 2875
rect 1025 2875 1075 2885
rect 1025 2855 1035 2875
rect 825 2850 1035 2855
rect 1065 2850 1075 2875
rect 425 2835 475 2850
rect 785 2840 1075 2850
rect 425 2810 435 2835
rect 465 2815 475 2835
rect 1385 2835 1435 2850
rect 1385 2815 1395 2835
rect 465 2810 1395 2815
rect 1425 2810 1435 2835
rect 425 2800 1435 2810
rect 920 2665 940 2800
rect 905 2655 955 2665
rect 360 2620 420 2640
rect 360 2600 380 2620
rect 400 2600 420 2620
rect -120 2580 -60 2595
rect 0 2580 60 2595
rect 120 2580 180 2595
rect 240 2580 300 2595
rect 360 2580 420 2600
rect 720 2620 780 2640
rect 905 2630 915 2655
rect 945 2630 955 2655
rect 905 2620 955 2630
rect 1080 2620 1140 2640
rect 1440 2635 1500 2655
rect 720 2600 740 2620
rect 760 2600 780 2620
rect 480 2580 540 2595
rect 600 2580 660 2595
rect 720 2580 780 2600
rect 1080 2600 1100 2620
rect 1120 2600 1140 2620
rect 840 2580 900 2595
rect 960 2580 1020 2595
rect 1080 2580 1140 2600
rect 1440 2615 1460 2635
rect 1480 2615 1500 2635
rect 1200 2580 1260 2595
rect 1320 2580 1380 2595
rect 1440 2580 1500 2615
rect 1560 2580 1620 2595
rect 1680 2580 1740 2595
rect 1800 2580 1860 2595
rect 1920 2580 1980 2595
rect -120 2415 -60 2430
rect -175 2405 -60 2415
rect -175 2385 -165 2405
rect -70 2385 -60 2405
rect -175 2375 -60 2385
rect 0 2390 60 2430
rect 120 2390 180 2430
rect 240 2390 300 2430
rect 360 2415 420 2430
rect 480 2390 540 2430
rect 600 2390 660 2430
rect 720 2415 780 2430
rect 840 2395 900 2430
rect 960 2395 1020 2430
rect 1080 2415 1140 2430
rect 840 2390 1020 2395
rect 1200 2390 1260 2430
rect 1320 2390 1380 2430
rect 1440 2415 1500 2430
rect 1560 2390 1620 2430
rect 1680 2390 1740 2430
rect 1800 2390 1860 2430
rect 0 2385 1860 2390
rect 0 2375 920 2385
rect 910 2365 920 2375
rect 940 2375 1860 2385
rect 1920 2415 1980 2430
rect 1920 2405 2035 2415
rect 1920 2385 1930 2405
rect 2025 2385 2035 2405
rect 1920 2375 2035 2385
rect 940 2365 950 2375
rect 910 2355 950 2365
<< polycont >>
rect 625 4850 645 4870
rect 1210 4850 1230 4870
rect -165 4630 -70 4650
rect -45 4630 50 4650
rect 75 4630 170 4650
rect 195 4630 290 4650
rect 315 4630 410 4650
rect 920 4560 940 4580
rect 1450 4630 1545 4650
rect 1570 4630 1665 4650
rect 1690 4630 1785 4650
rect 1810 4630 1905 4650
rect 1930 4630 2025 4650
rect 2030 4520 2050 4540
rect -165 4300 -70 4320
rect -45 4300 50 4320
rect 75 4300 170 4320
rect 195 4300 290 4320
rect 315 4300 410 4320
rect 735 4305 755 4325
rect 1105 4305 1125 4325
rect 1450 4300 1545 4320
rect 1570 4300 1665 4320
rect 1690 4300 1785 4320
rect 1810 4300 1905 4320
rect 1930 4300 2025 4320
rect -165 3855 -70 3875
rect -45 3855 50 3875
rect 75 3855 170 3875
rect 195 3855 290 3875
rect 490 3855 530 3875
rect 630 3855 650 3875
rect 850 3855 890 3875
rect 970 3855 1010 3875
rect 1210 3855 1230 3875
rect 1330 3855 1370 3875
rect 1570 3855 1665 3875
rect 1690 3855 1785 3875
rect 1810 3855 1905 3875
rect 1930 3855 2025 3875
rect 920 3795 940 3815
rect 920 3695 940 3715
rect 490 3635 530 3655
rect 630 3635 650 3655
rect 850 3635 890 3655
rect 970 3635 1010 3655
rect 1210 3635 1230 3655
rect 1330 3635 1370 3655
rect -165 3415 -70 3435
rect -45 3415 50 3435
rect 75 3415 170 3435
rect 195 3415 290 3435
rect 1570 3415 1665 3435
rect 1690 3415 1785 3435
rect 1810 3415 1905 3435
rect 1930 3415 2025 3435
rect 370 3160 390 3180
rect 440 3160 460 3180
rect 730 3160 750 3180
rect 1110 3160 1130 3180
rect 1470 3160 1490 3180
rect -165 2920 -70 2940
rect 1930 2920 2025 2940
rect 795 2850 825 2875
rect 1035 2850 1065 2875
rect 435 2810 465 2835
rect 1395 2810 1425 2835
rect 380 2600 400 2620
rect 915 2630 945 2655
rect 740 2600 760 2620
rect 1100 2600 1120 2620
rect 1460 2615 1480 2635
rect -165 2385 -70 2405
rect 920 2365 940 2385
rect 1930 2385 2025 2405
<< locali >>
rect 425 4950 1435 4970
rect 425 4915 475 4950
rect -225 4895 475 4915
rect -225 3330 -205 4895
rect -175 4810 -125 4820
rect -175 4690 -165 4810
rect -135 4690 -125 4810
rect -175 4660 -125 4690
rect -55 4810 -5 4820
rect -55 4690 -45 4810
rect -15 4690 -5 4810
rect -55 4660 -5 4690
rect 65 4810 115 4820
rect 65 4690 75 4810
rect 105 4690 115 4810
rect 65 4660 115 4690
rect 185 4810 235 4820
rect 185 4690 195 4810
rect 225 4690 235 4810
rect 185 4660 235 4690
rect 305 4810 355 4820
rect 305 4690 315 4810
rect 345 4690 355 4810
rect 305 4660 355 4690
rect 425 4810 475 4895
rect 425 4690 435 4810
rect 465 4690 475 4810
rect 425 4680 475 4690
rect 545 4910 1315 4930
rect 545 4810 595 4910
rect 615 4870 655 4880
rect 615 4850 625 4870
rect 645 4850 655 4870
rect 615 4840 655 4850
rect 545 4690 555 4810
rect 585 4690 595 4810
rect 545 4680 595 4690
rect 665 4810 715 4820
rect 665 4690 675 4810
rect 705 4690 715 4810
rect -175 4650 420 4660
rect -175 4630 -165 4650
rect -70 4630 -45 4650
rect 50 4630 75 4650
rect 170 4630 195 4650
rect 290 4630 315 4650
rect 410 4630 420 4650
rect -175 4620 420 4630
rect 665 4635 715 4690
rect 785 4810 835 4910
rect 785 4690 795 4810
rect 825 4690 835 4810
rect 785 4680 835 4690
rect 905 4810 955 4820
rect 905 4690 915 4810
rect 945 4690 955 4810
rect 905 4680 955 4690
rect 1025 4810 1075 4910
rect 1200 4870 1240 4880
rect 1200 4850 1210 4870
rect 1230 4850 1240 4870
rect 1200 4840 1240 4850
rect 1025 4690 1035 4810
rect 1065 4690 1075 4810
rect 1025 4680 1075 4690
rect 1145 4810 1195 4820
rect 1145 4690 1155 4810
rect 1185 4690 1195 4810
rect 1145 4635 1195 4690
rect 1265 4810 1315 4910
rect 1265 4690 1275 4810
rect 1305 4690 1315 4810
rect 1265 4680 1315 4690
rect 1385 4810 1435 4950
rect 1385 4690 1395 4810
rect 1425 4690 1435 4810
rect 1385 4680 1435 4690
rect 1505 4810 1555 4820
rect 1505 4690 1515 4810
rect 1545 4690 1555 4810
rect 1505 4660 1555 4690
rect 1625 4810 1675 4820
rect 1625 4690 1635 4810
rect 1665 4690 1675 4810
rect 1625 4660 1675 4690
rect 1745 4810 1795 4820
rect 1745 4690 1755 4810
rect 1785 4690 1795 4810
rect 1745 4660 1795 4690
rect 1865 4810 1915 4820
rect 1865 4690 1875 4810
rect 1905 4690 1915 4810
rect 1865 4660 1915 4690
rect 1985 4810 2035 4820
rect 1985 4690 1995 4810
rect 2025 4690 2035 4810
rect 1985 4660 2035 4690
rect 665 4615 1195 4635
rect 1440 4650 2035 4660
rect 1440 4630 1450 4650
rect 1545 4630 1570 4650
rect 1665 4630 1690 4650
rect 1785 4630 1810 4650
rect 1905 4630 1930 4650
rect 2025 4630 2035 4650
rect 1440 4620 2035 4630
rect 355 4595 405 4600
rect 170 4575 220 4585
rect 170 4545 180 4575
rect 210 4545 220 4575
rect 355 4565 365 4595
rect 395 4565 405 4595
rect 1465 4595 1515 4600
rect 355 4555 405 4565
rect 910 4580 950 4590
rect 910 4560 920 4580
rect 940 4570 950 4580
rect 940 4560 1235 4570
rect 910 4550 1235 4560
rect 1465 4565 1475 4595
rect 1505 4565 1515 4595
rect 1465 4555 1515 4565
rect 1725 4590 1775 4600
rect 1725 4560 1735 4590
rect 1765 4560 1775 4590
rect 1725 4550 1775 4560
rect 170 4535 220 4545
rect 1215 4530 1235 4550
rect 2020 4540 2060 4550
rect 2020 4530 2030 4540
rect 665 4510 1195 4530
rect 1215 4520 2030 4530
rect 2050 4520 2060 4540
rect 1215 4510 2060 4520
rect -175 4480 -125 4490
rect -175 4360 -165 4480
rect -135 4360 -125 4480
rect -175 4330 -125 4360
rect -55 4480 -5 4490
rect -55 4360 -45 4480
rect -15 4360 -5 4480
rect -55 4330 -5 4360
rect 65 4480 115 4490
rect 65 4360 75 4480
rect 105 4360 115 4480
rect 65 4330 115 4360
rect 185 4480 235 4490
rect 185 4360 195 4480
rect 225 4360 235 4480
rect 185 4330 235 4360
rect 305 4480 355 4490
rect 305 4360 315 4480
rect 345 4360 355 4480
rect 305 4330 355 4360
rect 425 4480 475 4490
rect 425 4360 435 4480
rect 465 4360 475 4480
rect 425 4350 475 4360
rect -175 4320 420 4330
rect -175 4300 -165 4320
rect -70 4300 -45 4320
rect 50 4300 75 4320
rect 170 4300 195 4320
rect 290 4300 315 4320
rect 410 4300 420 4320
rect -175 4290 420 4300
rect 455 4235 475 4350
rect 545 4480 595 4490
rect 545 4360 555 4480
rect 585 4360 595 4480
rect 545 4275 595 4360
rect 665 4480 715 4510
rect 665 4360 675 4480
rect 705 4360 715 4480
rect 665 4350 715 4360
rect 785 4480 835 4490
rect 785 4360 795 4480
rect 825 4360 835 4480
rect 725 4325 765 4335
rect 725 4305 735 4325
rect 755 4305 765 4325
rect 725 4295 765 4305
rect 785 4275 835 4360
rect 905 4480 955 4490
rect 905 4360 915 4480
rect 945 4360 955 4480
rect 905 4350 955 4360
rect 1025 4480 1075 4490
rect 1025 4360 1035 4480
rect 1065 4360 1075 4480
rect 1025 4275 1075 4360
rect 1145 4480 1195 4510
rect 1145 4360 1155 4480
rect 1185 4360 1195 4480
rect 1145 4350 1195 4360
rect 1265 4480 1315 4490
rect 1265 4360 1275 4480
rect 1305 4360 1315 4480
rect 1095 4325 1135 4335
rect 1095 4305 1105 4325
rect 1125 4305 1135 4325
rect 1095 4295 1135 4305
rect 1265 4275 1315 4360
rect 545 4255 1315 4275
rect 1385 4480 1435 4490
rect 1385 4360 1395 4480
rect 1425 4360 1435 4480
rect 1385 4350 1435 4360
rect 1505 4480 1555 4490
rect 1505 4360 1515 4480
rect 1545 4360 1555 4480
rect 1385 4235 1405 4350
rect 1505 4330 1555 4360
rect 1625 4480 1675 4490
rect 1625 4360 1635 4480
rect 1665 4360 1675 4480
rect 1625 4330 1675 4360
rect 1745 4480 1795 4490
rect 1745 4360 1755 4480
rect 1785 4360 1795 4480
rect 1745 4330 1795 4360
rect 1865 4480 1915 4490
rect 1865 4360 1875 4480
rect 1905 4360 1915 4480
rect 1865 4330 1915 4360
rect 1985 4480 2035 4490
rect 1985 4360 1995 4480
rect 2025 4360 2035 4480
rect 1985 4330 2035 4360
rect 1440 4320 2035 4330
rect 1440 4300 1450 4320
rect 1545 4300 1570 4320
rect 1665 4300 1690 4320
rect 1785 4300 1810 4320
rect 1905 4300 1930 4320
rect 2025 4300 2035 4320
rect 1440 4290 2035 4300
rect 455 4215 1405 4235
rect 455 4195 475 4215
rect 1385 4195 1405 4215
rect 455 4175 2080 4195
rect 455 4050 475 4175
rect -175 4035 -125 4045
rect -175 3915 -165 4035
rect -135 3915 -125 4035
rect -175 3885 -125 3915
rect -55 4035 -5 4045
rect -55 3915 -45 4035
rect -15 3915 -5 4035
rect -55 3885 -5 3915
rect 65 4035 115 4045
rect 65 3915 75 4035
rect 105 3915 115 4035
rect 65 3885 115 3915
rect 185 4035 235 4045
rect 185 3915 195 4035
rect 225 3915 235 4035
rect 185 3885 235 3915
rect 305 4035 355 4045
rect 305 3915 315 4035
rect 345 3915 355 4035
rect 305 3905 355 3915
rect 425 4035 475 4050
rect 785 4135 1075 4155
rect 425 3915 435 4035
rect 465 3915 475 4035
rect 425 3905 475 3915
rect 545 4035 595 4045
rect 545 3915 555 4035
rect 585 3915 595 4035
rect 545 3885 595 3915
rect 665 4035 715 4045
rect 665 3915 675 4035
rect 705 3915 715 4035
rect 665 3885 715 3915
rect 785 4035 835 4135
rect 785 3915 795 4035
rect 825 3915 835 4035
rect 785 3905 835 3915
rect 905 4035 955 4045
rect 905 3915 915 4035
rect 945 3915 955 4035
rect 905 3905 955 3915
rect 1025 4035 1075 4135
rect 1385 4050 1405 4175
rect 1025 3915 1035 4035
rect 1065 3915 1075 4035
rect 1025 3905 1075 3915
rect 1145 4035 1195 4045
rect 1145 3915 1155 4035
rect 1185 3915 1195 4035
rect -175 3875 300 3885
rect -175 3855 -165 3875
rect -70 3855 -45 3875
rect 50 3855 75 3875
rect 170 3855 195 3875
rect 290 3855 300 3875
rect -175 3845 300 3855
rect 480 3875 595 3885
rect 480 3855 490 3875
rect 530 3855 595 3875
rect 480 3845 595 3855
rect 620 3875 715 3885
rect 620 3855 630 3875
rect 650 3865 715 3875
rect 840 3875 900 3885
rect 650 3855 660 3865
rect 620 3845 660 3855
rect 840 3855 850 3875
rect 890 3855 900 3875
rect 840 3845 900 3855
rect 365 3835 415 3845
rect 365 3800 375 3835
rect 405 3800 415 3835
rect 365 3790 415 3800
rect 480 3765 540 3845
rect 840 3765 890 3845
rect 920 3825 940 3905
rect 1145 3885 1195 3915
rect 1265 4035 1315 4045
rect 1265 3915 1275 4035
rect 1305 3915 1315 4035
rect 1265 3885 1315 3915
rect 1385 4035 1435 4050
rect 1385 3915 1395 4035
rect 1425 3915 1435 4035
rect 1385 3905 1435 3915
rect 1505 4035 1555 4045
rect 1505 3915 1515 4035
rect 1545 3915 1555 4035
rect 1505 3905 1555 3915
rect 1625 4035 1675 4045
rect 1625 3915 1635 4035
rect 1665 3915 1675 4035
rect 1625 3885 1675 3915
rect 1745 4035 1795 4045
rect 1745 3915 1755 4035
rect 1785 3915 1795 4035
rect 1745 3885 1795 3915
rect 1865 4035 1915 4045
rect 1865 3915 1875 4035
rect 1905 3915 1915 4035
rect 1865 3885 1915 3915
rect 1985 4035 2035 4045
rect 1985 3915 1995 4035
rect 2025 3915 2035 4035
rect 1985 3885 2035 3915
rect 960 3875 1020 3885
rect 960 3855 970 3875
rect 1010 3855 1020 3875
rect 1145 3875 1240 3885
rect 1145 3865 1210 3875
rect 960 3845 1020 3855
rect 1200 3855 1210 3865
rect 1230 3855 1240 3875
rect 1200 3845 1240 3855
rect 1265 3875 1380 3885
rect 1265 3855 1330 3875
rect 1370 3855 1380 3875
rect 1265 3845 1380 3855
rect 1560 3875 2035 3885
rect 1560 3855 1570 3875
rect 1665 3855 1690 3875
rect 1785 3855 1810 3875
rect 1905 3855 1930 3875
rect 2025 3855 2035 3875
rect 1560 3845 2035 3855
rect 910 3815 950 3825
rect 910 3795 920 3815
rect 940 3795 950 3815
rect 910 3785 950 3795
rect 970 3765 1020 3845
rect 1320 3765 1380 3845
rect 1445 3825 1495 3835
rect 1445 3790 1455 3825
rect 1485 3790 1495 3825
rect 1445 3780 1495 3790
rect 170 3755 220 3765
rect 170 3720 180 3755
rect 210 3720 220 3755
rect 170 3710 220 3720
rect 480 3745 1380 3765
rect 480 3665 540 3745
rect 840 3665 890 3745
rect 910 3715 950 3725
rect 910 3695 920 3715
rect 940 3695 950 3715
rect 910 3685 950 3695
rect 480 3655 595 3665
rect 480 3635 490 3655
rect 530 3635 595 3655
rect 480 3625 595 3635
rect 620 3655 660 3665
rect 620 3635 630 3655
rect 650 3645 660 3655
rect 840 3655 900 3665
rect 650 3635 715 3645
rect 620 3625 715 3635
rect 840 3635 850 3655
rect 890 3635 900 3655
rect 840 3625 900 3635
rect -175 3595 -125 3605
rect -175 3475 -165 3595
rect -135 3475 -125 3595
rect -175 3445 -125 3475
rect -55 3595 -5 3605
rect -55 3475 -45 3595
rect -15 3475 -5 3595
rect -55 3445 -5 3475
rect 65 3595 115 3605
rect 65 3475 75 3595
rect 105 3475 115 3595
rect 65 3445 115 3475
rect 185 3595 235 3605
rect 185 3475 195 3595
rect 225 3475 235 3595
rect 185 3445 235 3475
rect 305 3595 355 3605
rect 305 3475 315 3595
rect 345 3475 355 3595
rect 305 3465 355 3475
rect 425 3595 475 3605
rect 425 3475 435 3595
rect 465 3475 475 3595
rect -175 3435 300 3445
rect -175 3415 -165 3435
rect -70 3415 -45 3435
rect 50 3415 75 3435
rect 170 3415 195 3435
rect 290 3415 300 3435
rect -175 3405 300 3415
rect 425 3330 475 3475
rect 545 3595 595 3625
rect 545 3475 555 3595
rect 585 3475 595 3595
rect 545 3465 595 3475
rect 665 3595 715 3625
rect 920 3605 940 3685
rect 970 3665 1020 3745
rect 1320 3665 1380 3745
rect 1680 3745 1730 3755
rect 1680 3710 1690 3745
rect 1720 3710 1730 3745
rect 1680 3700 1730 3710
rect 960 3655 1020 3665
rect 960 3635 970 3655
rect 1010 3635 1020 3655
rect 1200 3655 1240 3665
rect 1200 3645 1210 3655
rect 960 3625 1020 3635
rect 1145 3635 1210 3645
rect 1230 3635 1240 3655
rect 1145 3625 1240 3635
rect 1265 3655 1380 3665
rect 1265 3635 1330 3655
rect 1370 3635 1380 3655
rect 1265 3625 1380 3635
rect 665 3475 675 3595
rect 705 3475 715 3595
rect 665 3465 715 3475
rect 785 3595 835 3605
rect 785 3475 795 3595
rect 825 3475 835 3595
rect 785 3370 835 3475
rect 905 3595 955 3605
rect 905 3475 915 3595
rect 945 3475 955 3595
rect 905 3465 955 3475
rect 1025 3595 1075 3605
rect 1025 3475 1035 3595
rect 1065 3475 1075 3595
rect 1025 3370 1075 3475
rect 1145 3595 1195 3625
rect 1145 3475 1155 3595
rect 1185 3475 1195 3595
rect 1145 3465 1195 3475
rect 1265 3595 1315 3625
rect 1265 3475 1275 3595
rect 1305 3475 1315 3595
rect 1265 3465 1315 3475
rect 1385 3595 1435 3605
rect 1385 3475 1395 3595
rect 1425 3475 1435 3595
rect 785 3350 1075 3370
rect 1385 3330 1435 3475
rect 1505 3595 1555 3605
rect 1505 3475 1515 3595
rect 1545 3475 1555 3595
rect 1505 3465 1555 3475
rect 1625 3595 1675 3605
rect 1625 3475 1635 3595
rect 1665 3475 1675 3595
rect 1625 3445 1675 3475
rect 1745 3595 1795 3605
rect 1745 3475 1755 3595
rect 1785 3475 1795 3595
rect 1745 3445 1795 3475
rect 1865 3595 1915 3605
rect 1865 3475 1875 3595
rect 1905 3475 1915 3595
rect 1865 3445 1915 3475
rect 1985 3595 2035 3605
rect 1985 3475 1995 3595
rect 2025 3475 2035 3595
rect 1985 3445 2035 3475
rect 1560 3435 2035 3445
rect 1560 3415 1570 3435
rect 1665 3415 1690 3435
rect 1785 3415 1810 3435
rect 1905 3415 1930 3435
rect 2025 3415 2035 3435
rect 1560 3405 2035 3415
rect -225 3320 1435 3330
rect -225 3310 920 3320
rect 910 3300 920 3310
rect 940 3310 1435 3320
rect 940 3300 950 3310
rect 910 3290 950 3300
rect 2060 3290 2080 4175
rect 1030 3280 2080 3290
rect 1030 3260 1040 3280
rect 1060 3260 2080 3280
rect 1030 3250 2080 3260
rect 65 3210 1795 3230
rect -175 3100 -125 3110
rect -175 2980 -165 3100
rect -135 2980 -125 3100
rect -175 2950 -125 2980
rect -55 3100 -5 3110
rect -55 2980 -45 3100
rect -15 2980 -5 3100
rect -55 2970 -5 2980
rect 65 3100 115 3210
rect 305 3115 325 3210
rect 360 3180 400 3190
rect 360 3160 370 3180
rect 390 3160 400 3180
rect 360 3150 400 3160
rect 430 3180 470 3190
rect 430 3160 440 3180
rect 460 3160 470 3180
rect 430 3150 470 3160
rect 65 2980 75 3100
rect 105 2980 115 3100
rect 65 2970 115 2980
rect 185 3100 235 3110
rect 185 2980 195 3100
rect 225 2980 235 3100
rect 185 2970 235 2980
rect 305 3100 355 3115
rect 305 2980 315 3100
rect 345 2980 355 3100
rect 305 2970 355 2980
rect 425 3100 475 3150
rect 425 2980 435 3100
rect 465 2980 475 3100
rect -175 2940 -60 2950
rect -175 2920 -165 2940
rect -70 2920 -60 2940
rect -175 2910 -60 2920
rect 240 2870 350 2880
rect 240 2780 250 2870
rect 340 2780 350 2870
rect 425 2835 475 2980
rect 545 3100 595 3210
rect 720 3180 760 3190
rect 720 3160 730 3180
rect 750 3160 760 3180
rect 720 3150 760 3160
rect 1100 3180 1140 3190
rect 1100 3160 1110 3180
rect 1130 3160 1140 3180
rect 1100 3150 1140 3160
rect 545 2980 555 3100
rect 585 2980 595 3100
rect 545 2970 595 2980
rect 665 3100 715 3110
rect 665 2980 675 3100
rect 705 2980 715 3100
rect 665 2970 715 2980
rect 785 3100 835 3110
rect 785 2980 795 3100
rect 825 2980 835 3100
rect 785 2875 835 2980
rect 785 2850 795 2875
rect 825 2850 835 2875
rect 785 2840 835 2850
rect 905 3100 955 3110
rect 905 2980 915 3100
rect 945 2980 955 3100
rect 425 2810 435 2835
rect 465 2810 475 2835
rect 425 2800 475 2810
rect 240 2770 350 2780
rect 905 2755 955 2980
rect 1025 3100 1075 3110
rect 1025 2980 1035 3100
rect 1065 2980 1075 3100
rect 1025 2875 1075 2980
rect 1145 3100 1195 3110
rect 1145 2980 1155 3100
rect 1185 2980 1195 3100
rect 1145 2970 1195 2980
rect 1265 3100 1315 3210
rect 1460 3180 1500 3190
rect 1460 3160 1470 3180
rect 1490 3160 1500 3180
rect 1460 3150 1500 3160
rect 1535 3115 1555 3210
rect 1265 2980 1275 3100
rect 1305 2980 1315 3100
rect 1265 2970 1315 2980
rect 1385 3100 1435 3110
rect 1385 2980 1395 3100
rect 1425 2980 1435 3100
rect 1025 2850 1035 2875
rect 1065 2850 1075 2875
rect 1025 2840 1075 2850
rect 1385 2835 1435 2980
rect 1505 3100 1555 3115
rect 1505 2980 1515 3100
rect 1545 2980 1555 3100
rect 1505 2970 1555 2980
rect 1625 3100 1675 3110
rect 1625 2980 1635 3100
rect 1665 2980 1675 3100
rect 1625 2970 1675 2980
rect 1745 3100 1795 3210
rect 1745 2980 1755 3100
rect 1785 2980 1795 3100
rect 1745 2970 1795 2980
rect 1865 3100 1915 3110
rect 1865 2980 1875 3100
rect 1905 2980 1915 3100
rect 1865 2970 1915 2980
rect 1985 3100 2035 3110
rect 1985 2980 1995 3100
rect 2025 2980 2035 3100
rect 1985 2950 2035 2980
rect 1920 2940 2035 2950
rect 1920 2920 1930 2940
rect 2025 2920 2035 2940
rect 1920 2910 2035 2920
rect 1385 2810 1395 2835
rect 1425 2810 1435 2835
rect 1385 2800 1435 2810
rect 1520 2870 1630 2880
rect 1520 2780 1530 2870
rect 1620 2780 1630 2870
rect 1520 2770 1630 2780
rect 455 2730 565 2740
rect 455 2640 465 2730
rect 555 2640 565 2730
rect 455 2630 565 2640
rect 665 2735 1195 2755
rect 370 2620 410 2630
rect 370 2600 380 2620
rect 400 2600 410 2620
rect 370 2590 410 2600
rect 665 2580 685 2735
rect 815 2695 920 2705
rect 940 2695 1045 2705
rect 815 2685 1045 2695
rect 730 2620 770 2630
rect 730 2600 740 2620
rect 760 2600 770 2620
rect 730 2590 770 2600
rect 815 2580 835 2685
rect -175 2565 -125 2575
rect -175 2445 -165 2565
rect -135 2445 -125 2565
rect -175 2415 -125 2445
rect -55 2565 -5 2575
rect -55 2445 -45 2565
rect -15 2445 -5 2565
rect -55 2435 -5 2445
rect 65 2565 115 2575
rect 65 2445 75 2565
rect 105 2445 115 2565
rect -175 2405 -60 2415
rect -175 2385 -165 2405
rect -70 2385 -60 2405
rect -175 2375 -60 2385
rect 65 2335 115 2445
rect 185 2565 235 2575
rect 185 2445 195 2565
rect 225 2445 235 2565
rect 185 2435 235 2445
rect 305 2565 355 2575
rect 305 2445 315 2565
rect 345 2445 355 2565
rect 305 2335 355 2445
rect 425 2565 475 2575
rect 425 2445 435 2565
rect 465 2445 475 2565
rect 425 2435 475 2445
rect 545 2565 595 2575
rect 545 2445 555 2565
rect 585 2445 595 2565
rect 545 2335 595 2445
rect 665 2565 715 2580
rect 665 2445 675 2565
rect 705 2445 715 2565
rect 665 2435 715 2445
rect 785 2565 835 2580
rect 785 2445 795 2565
rect 825 2445 835 2565
rect 785 2435 835 2445
rect 905 2655 955 2665
rect 905 2630 915 2655
rect 945 2630 955 2655
rect 905 2565 955 2630
rect 905 2445 915 2565
rect 945 2445 955 2565
rect 905 2435 955 2445
rect 1025 2580 1045 2685
rect 1090 2620 1130 2630
rect 1090 2600 1100 2620
rect 1120 2600 1130 2620
rect 1090 2590 1130 2600
rect 1175 2580 1195 2735
rect 1295 2730 1405 2740
rect 1295 2640 1305 2730
rect 1395 2640 1405 2730
rect 1295 2630 1405 2640
rect 1450 2635 1490 2645
rect 1450 2615 1460 2635
rect 1480 2615 1490 2635
rect 1450 2605 1490 2615
rect 1025 2565 1075 2580
rect 1025 2445 1035 2565
rect 1065 2445 1075 2565
rect 1025 2435 1075 2445
rect 1145 2565 1195 2580
rect 1145 2445 1155 2565
rect 1185 2445 1195 2565
rect 1145 2435 1195 2445
rect 1265 2565 1315 2575
rect 1265 2445 1275 2565
rect 1305 2445 1315 2565
rect 910 2385 950 2435
rect 910 2365 920 2385
rect 940 2365 950 2385
rect 910 2355 950 2365
rect 1265 2335 1315 2445
rect 1385 2565 1435 2575
rect 1385 2445 1395 2565
rect 1425 2445 1435 2565
rect 1385 2435 1435 2445
rect 1505 2565 1555 2575
rect 1505 2445 1515 2565
rect 1545 2445 1555 2565
rect 1505 2335 1555 2445
rect 1625 2565 1675 2575
rect 1625 2445 1635 2565
rect 1665 2445 1675 2565
rect 1625 2435 1675 2445
rect 1745 2565 1795 2575
rect 1745 2445 1755 2565
rect 1785 2445 1795 2565
rect 1745 2335 1795 2445
rect 1865 2565 1915 2575
rect 1865 2445 1875 2565
rect 1905 2445 1915 2565
rect 1865 2435 1915 2445
rect 1985 2565 2035 2575
rect 1985 2445 1995 2565
rect 2025 2445 2035 2565
rect 1985 2415 2035 2445
rect 1920 2405 2035 2415
rect 1920 2385 1930 2405
rect 2025 2385 2035 2405
rect 1920 2375 2035 2385
rect 65 2315 1795 2335
<< viali >>
rect -165 4690 -135 4810
rect -45 4690 -15 4810
rect 75 4690 105 4810
rect 195 4690 225 4810
rect 315 4690 345 4810
rect 915 4690 945 4810
rect 1515 4690 1545 4810
rect 1635 4690 1665 4810
rect 1755 4690 1785 4810
rect 1875 4690 1905 4810
rect 1995 4690 2025 4810
rect 180 4545 210 4575
rect 365 4565 395 4595
rect 1475 4565 1505 4595
rect 1735 4560 1765 4590
rect -165 4360 -135 4480
rect -45 4360 -15 4480
rect 75 4360 105 4480
rect 195 4360 225 4480
rect 315 4360 345 4480
rect 735 4305 755 4325
rect 915 4360 945 4480
rect 1105 4305 1125 4325
rect 1515 4360 1545 4480
rect 1635 4360 1665 4480
rect 1755 4360 1785 4480
rect 1875 4360 1905 4480
rect 1995 4360 2025 4480
rect -165 3915 -135 4035
rect -45 3915 -15 4035
rect 75 3915 105 4035
rect 195 3915 225 4035
rect 315 3915 345 4035
rect 675 3915 705 4035
rect 1155 3915 1185 4035
rect 375 3800 405 3835
rect 1515 3915 1545 4035
rect 1635 3915 1665 4035
rect 1755 3915 1785 4035
rect 1875 3915 1905 4035
rect 1995 3915 2025 4035
rect 1455 3790 1485 3825
rect 180 3720 210 3755
rect -165 3475 -135 3595
rect -45 3475 -15 3595
rect 75 3475 105 3595
rect 195 3475 225 3595
rect 315 3475 345 3595
rect 1690 3710 1720 3745
rect 675 3475 705 3595
rect 1155 3475 1185 3595
rect 1515 3475 1545 3595
rect 1635 3475 1665 3595
rect 1755 3475 1785 3595
rect 1875 3475 1905 3595
rect 1995 3475 2025 3595
rect 920 3300 940 3320
rect 1040 3260 1060 3280
rect -165 2980 -135 3100
rect -45 2980 -15 3100
rect 370 3160 390 3180
rect 195 2980 225 3100
rect 250 2780 340 2870
rect 730 3160 750 3180
rect 1110 3160 1130 3180
rect 675 2980 705 3100
rect 1155 2980 1185 3100
rect 1470 3160 1490 3180
rect 1035 2850 1065 2875
rect 1635 2980 1665 3100
rect 1875 2980 1905 3100
rect 1995 2980 2025 3100
rect 1530 2780 1620 2870
rect 465 2640 555 2730
rect 380 2600 400 2620
rect 920 2695 940 2715
rect 740 2600 760 2620
rect -165 2445 -135 2565
rect -45 2445 -15 2565
rect 195 2445 225 2565
rect 435 2445 465 2565
rect 1100 2600 1120 2620
rect 1305 2640 1395 2730
rect 1460 2615 1480 2635
rect 1395 2445 1425 2565
rect 1635 2445 1665 2565
rect 1875 2445 1905 2565
rect 1995 2445 2025 2565
<< metal1 >>
rect -250 4810 595 4820
rect -250 4690 -165 4810
rect -135 4690 -45 4810
rect -15 4690 75 4810
rect 105 4690 195 4810
rect 225 4690 315 4810
rect 345 4690 595 4810
rect -250 4680 595 4690
rect 905 4810 955 4820
rect 905 4690 915 4810
rect 945 4690 955 4810
rect 905 4680 955 4690
rect 1265 4810 2110 4820
rect 1265 4690 1515 4810
rect 1545 4690 1635 4810
rect 1665 4690 1755 4810
rect 1785 4690 1875 4810
rect 1905 4690 1995 4810
rect 2025 4690 2110 4810
rect 1265 4680 2110 4690
rect -250 4045 -200 4680
rect 165 4575 225 4680
rect 165 4545 180 4575
rect 210 4545 225 4575
rect 350 4595 410 4605
rect 350 4565 365 4595
rect 395 4565 410 4595
rect 350 4550 410 4565
rect 165 4530 225 4545
rect 545 4490 595 4680
rect 1265 4490 1315 4680
rect 1460 4595 1520 4605
rect 1460 4565 1475 4595
rect 1505 4565 1520 4595
rect 1460 4550 1520 4565
rect 1720 4590 1780 4680
rect 1720 4560 1735 4590
rect 1765 4560 1780 4590
rect 1720 4545 1780 4560
rect -175 4480 -125 4490
rect -175 4360 -165 4480
rect -135 4360 -125 4480
rect -175 4350 -125 4360
rect -55 4480 -5 4490
rect -55 4360 -45 4480
rect -15 4360 -5 4480
rect -55 4350 -5 4360
rect 65 4480 115 4490
rect 65 4360 75 4480
rect 105 4360 115 4480
rect 65 4350 115 4360
rect 185 4480 235 4490
rect 185 4360 195 4480
rect 225 4360 235 4480
rect 185 4350 235 4360
rect 305 4480 355 4490
rect 305 4360 315 4480
rect 345 4360 355 4480
rect 305 4350 355 4360
rect 545 4480 1315 4490
rect 545 4360 915 4480
rect 945 4360 1315 4480
rect 545 4350 1315 4360
rect 1505 4480 1555 4490
rect 1505 4360 1515 4480
rect 1545 4360 1555 4480
rect 1505 4350 1555 4360
rect 1625 4480 1675 4490
rect 1625 4360 1635 4480
rect 1665 4360 1675 4480
rect 1625 4350 1675 4360
rect 1745 4480 1795 4490
rect 1745 4360 1755 4480
rect 1785 4360 1795 4480
rect 1745 4350 1795 4360
rect 1865 4480 1915 4490
rect 1865 4360 1875 4480
rect 1905 4360 1915 4480
rect 1865 4350 1915 4360
rect 1985 4480 2035 4490
rect 1985 4360 1995 4480
rect 2025 4360 2035 4480
rect 1985 4350 2035 4360
rect 720 4325 780 4350
rect 720 4305 735 4325
rect 755 4305 780 4325
rect 720 4295 780 4305
rect 1080 4325 1140 4350
rect 1080 4305 1105 4325
rect 1125 4305 1140 4325
rect 1080 4295 1140 4305
rect 2060 4045 2110 4680
rect -250 4035 240 4045
rect -250 3915 -165 4035
rect -135 3915 -45 4035
rect -15 3915 75 4035
rect 105 3915 195 4035
rect 225 3915 240 4035
rect -250 3905 240 3915
rect 305 4035 355 4045
rect 305 3915 315 4035
rect 345 3915 355 4035
rect 305 3905 355 3915
rect 665 4035 715 4045
rect 665 3915 675 4035
rect 705 3915 715 4035
rect 665 3905 715 3915
rect 1145 4035 1195 4045
rect 1145 3915 1155 4035
rect 1185 3915 1195 4035
rect 1145 3905 1195 3915
rect 1505 4035 1555 4045
rect 1505 3915 1515 4035
rect 1545 3915 1555 4035
rect 1505 3905 1555 3915
rect 1625 4035 2110 4045
rect 1625 3915 1635 4035
rect 1665 3915 1755 4035
rect 1785 3915 1875 4035
rect 1905 3915 1995 4035
rect 2025 3915 2110 4035
rect 1625 3905 2110 3915
rect 165 3900 240 3905
rect 165 3755 225 3900
rect 365 3835 415 3845
rect 365 3800 375 3835
rect 405 3800 415 3835
rect 365 3790 415 3800
rect 1445 3825 1495 3835
rect 1445 3790 1455 3825
rect 1485 3790 1495 3825
rect 1445 3780 1495 3790
rect 165 3720 180 3755
rect 210 3720 225 3755
rect 165 3685 225 3720
rect 1675 3745 1735 3905
rect 1675 3710 1690 3745
rect 1720 3710 1735 3745
rect 1675 3685 1735 3710
rect 165 3635 355 3685
rect 305 3605 355 3635
rect 1505 3635 1735 3685
rect 1505 3605 1555 3635
rect -175 3595 -125 3605
rect -175 3475 -165 3595
rect -135 3475 -125 3595
rect -175 3465 -125 3475
rect -55 3595 -5 3605
rect -55 3475 -45 3595
rect -15 3475 -5 3595
rect -55 3465 -5 3475
rect 65 3595 115 3605
rect 65 3475 75 3595
rect 105 3475 115 3595
rect 65 3465 115 3475
rect 185 3595 235 3605
rect 185 3475 195 3595
rect 225 3475 235 3595
rect 185 3465 235 3475
rect 305 3595 715 3605
rect 305 3475 315 3595
rect 345 3475 675 3595
rect 705 3475 715 3595
rect 305 3465 715 3475
rect 1145 3595 1555 3605
rect 1145 3475 1155 3595
rect 1185 3475 1515 3595
rect 1545 3475 1555 3595
rect 1145 3465 1555 3475
rect 1625 3595 1675 3605
rect 1625 3475 1635 3595
rect 1665 3475 1675 3595
rect 1625 3465 1675 3475
rect 1745 3595 1795 3605
rect 1745 3475 1755 3595
rect 1785 3475 1795 3595
rect 1745 3465 1795 3475
rect 1865 3595 1915 3605
rect 1865 3475 1875 3595
rect 1905 3475 1915 3595
rect 1865 3465 1915 3475
rect 1985 3595 2035 3605
rect 1985 3475 1995 3595
rect 2025 3475 2035 3595
rect 1985 3465 2035 3475
rect 305 3260 355 3465
rect 180 3210 355 3260
rect 910 3320 950 3330
rect 910 3300 920 3320
rect 940 3300 950 3320
rect -180 3110 -120 3115
rect 180 3110 235 3210
rect -180 3100 235 3110
rect -180 2980 -165 3100
rect -135 2980 -45 3100
rect -15 2980 195 3100
rect 225 2980 235 3100
rect -180 2970 235 2980
rect 355 3180 405 3190
rect 355 3160 370 3180
rect 390 3160 405 3180
rect 355 3110 405 3160
rect 720 3180 765 3190
rect 720 3160 730 3180
rect 750 3160 765 3180
rect 720 3110 765 3160
rect 355 3100 785 3110
rect 355 2980 675 3100
rect 705 2980 785 3100
rect 355 2970 785 2980
rect -180 2690 -5 2970
rect 355 2885 405 2970
rect 235 2870 405 2885
rect 235 2780 250 2870
rect 340 2780 405 2870
rect 235 2765 405 2780
rect 420 2730 600 2755
rect 420 2690 465 2730
rect -180 2640 465 2690
rect 555 2640 600 2730
rect 910 2715 950 3300
rect 1025 3280 1075 3295
rect 1025 3260 1040 3280
rect 1060 3260 1075 3280
rect 1025 2875 1075 3260
rect 1505 3260 1555 3465
rect 1505 3210 1675 3260
rect 1095 3180 1140 3190
rect 1095 3160 1110 3180
rect 1130 3160 1140 3180
rect 1095 3110 1140 3160
rect 1450 3180 1500 3190
rect 1450 3160 1470 3180
rect 1490 3160 1500 3180
rect 1450 3110 1500 3160
rect 1095 3100 1500 3110
rect 1095 2980 1155 3100
rect 1185 2980 1500 3100
rect 1095 2970 1500 2980
rect 1625 3110 1675 3210
rect 1625 3100 2040 3110
rect 1625 2980 1635 3100
rect 1665 2980 1875 3100
rect 1905 2980 1995 3100
rect 2025 2980 2040 3100
rect 1625 2970 2040 2980
rect 1025 2850 1035 2875
rect 1065 2850 1075 2875
rect 1025 2840 1075 2850
rect 1450 2885 1500 2970
rect 1450 2870 1635 2885
rect 1450 2780 1530 2870
rect 1620 2780 1635 2870
rect 1450 2765 1635 2780
rect 910 2695 920 2715
rect 940 2695 950 2715
rect 910 2685 950 2695
rect 1260 2730 1440 2755
rect 1260 2640 1305 2730
rect 1395 2705 1440 2730
rect 1865 2705 2035 2970
rect 1395 2655 2035 2705
rect 1395 2640 1500 2655
rect 360 2620 600 2640
rect 360 2600 380 2620
rect 400 2600 600 2620
rect 360 2580 600 2600
rect 720 2620 780 2640
rect 720 2600 740 2620
rect 760 2600 780 2620
rect 720 2580 780 2600
rect 1080 2620 1140 2640
rect 1080 2600 1100 2620
rect 1120 2600 1140 2620
rect 1080 2580 1140 2600
rect 1260 2635 1500 2640
rect 1260 2615 1460 2635
rect 1480 2615 1500 2635
rect 1260 2580 1500 2615
rect -175 2565 -125 2575
rect -175 2445 -165 2565
rect -135 2445 -125 2565
rect -175 2435 -125 2445
rect -55 2565 -5 2575
rect -55 2445 -45 2565
rect -15 2445 -5 2565
rect -55 2435 -5 2445
rect 185 2565 235 2575
rect 185 2445 195 2565
rect 225 2445 235 2565
rect 185 2435 235 2445
rect 360 2565 1500 2580
rect 360 2445 435 2565
rect 465 2445 1395 2565
rect 1425 2445 1500 2565
rect 360 2430 1500 2445
rect 1625 2565 1675 2575
rect 1625 2445 1635 2565
rect 1665 2445 1675 2565
rect 1625 2435 1675 2445
rect 1865 2565 1915 2575
rect 1865 2445 1875 2565
rect 1905 2445 1915 2565
rect 1865 2435 1915 2445
rect 1985 2565 2035 2575
rect 1985 2445 1995 2565
rect 2025 2445 2035 2565
rect 1985 2435 2035 2445
<< via1 >>
rect 915 4690 945 4810
rect 365 4565 395 4595
rect 1475 4565 1505 4595
rect -165 4360 -135 4480
rect -45 4360 -15 4480
rect 75 4360 105 4480
rect 195 4360 225 4480
rect 315 4360 345 4480
rect 1515 4360 1545 4480
rect 1635 4360 1665 4480
rect 1755 4360 1785 4480
rect 1875 4360 1905 4480
rect 1995 4360 2025 4480
rect 315 3915 345 4035
rect 675 3915 705 4035
rect 1155 3915 1185 4035
rect 1515 3915 1545 4035
rect 375 3800 405 3835
rect 1455 3790 1485 3825
rect -165 3475 -135 3595
rect -45 3475 -15 3595
rect 75 3475 105 3595
rect 195 3475 225 3595
rect 1635 3475 1665 3595
rect 1755 3475 1785 3595
rect 1875 3475 1905 3595
rect 1995 3475 2025 3595
rect 250 2780 340 2870
rect 1530 2780 1620 2870
rect -165 2445 -135 2565
rect -45 2445 -15 2565
rect 195 2445 225 2565
rect 1635 2445 1665 2565
rect 1875 2445 1905 2565
rect 1995 2445 2025 2565
<< metal2 >>
rect 605 4605 655 4880
rect 905 4810 955 4820
rect 905 4690 915 4810
rect 945 4690 955 4810
rect 905 4605 955 4690
rect 1200 4605 1260 4880
rect 305 4595 1555 4605
rect 305 4565 365 4595
rect 395 4565 1475 4595
rect 1505 4565 1555 4595
rect 305 4555 1555 4565
rect 305 4550 410 4555
rect 1460 4550 1555 4555
rect 305 4490 355 4550
rect -180 4480 355 4490
rect -180 4360 -165 4480
rect -135 4360 -45 4480
rect -15 4360 75 4480
rect 105 4360 195 4480
rect 225 4360 315 4480
rect 345 4360 355 4480
rect -180 4350 355 4360
rect 305 4045 355 4350
rect 1505 4490 1555 4550
rect 1505 4480 2035 4490
rect 1505 4360 1515 4480
rect 1545 4360 1635 4480
rect 1665 4360 1755 4480
rect 1785 4360 1875 4480
rect 1905 4360 1995 4480
rect 2025 4360 2035 4480
rect 1505 4350 2035 4360
rect 1505 4045 1555 4350
rect 305 4035 715 4045
rect 305 3915 315 4035
rect 345 3915 675 4035
rect 705 3915 715 4035
rect 305 3905 715 3915
rect 1145 4035 1555 4045
rect 1145 3915 1155 4035
rect 1185 3915 1515 4035
rect 1545 3915 1555 4035
rect 1145 3905 1555 3915
rect 355 3835 425 3905
rect 355 3800 375 3835
rect 405 3800 425 3835
rect 355 3605 425 3800
rect 1445 3825 1495 3905
rect 1445 3790 1455 3825
rect 1485 3790 1495 3825
rect 1445 3605 1495 3790
rect -180 3595 435 3605
rect -180 3475 -165 3595
rect -135 3475 -45 3595
rect -15 3475 75 3595
rect 105 3475 195 3595
rect 225 3475 435 3595
rect -180 3465 435 3475
rect 1445 3595 2035 3605
rect 1445 3475 1635 3595
rect 1665 3475 1755 3595
rect 1785 3475 1875 3595
rect 1905 3475 1995 3595
rect 2025 3475 2035 3595
rect 1445 3465 2035 3475
rect -175 2575 -5 3465
rect 355 3460 425 3465
rect 180 2870 355 2885
rect 180 2780 250 2870
rect 340 2780 355 2870
rect 180 2765 355 2780
rect 1515 2870 1675 2885
rect 1515 2780 1530 2870
rect 1620 2780 1675 2870
rect 1515 2765 1675 2780
rect 180 2575 240 2765
rect -180 2565 240 2575
rect -180 2445 -165 2565
rect -135 2445 -45 2565
rect -15 2445 195 2565
rect 225 2445 240 2565
rect -180 2435 240 2445
rect 1625 2575 1675 2765
rect 1865 2575 2035 3465
rect 1625 2565 2040 2575
rect 1625 2445 1635 2565
rect 1665 2445 1875 2565
rect 1905 2445 1995 2565
rect 2025 2445 2040 2565
rect 1625 2435 2040 2445
<< end >>
