magic
tech sky130A
timestamp 1620758016
<< locali >>
rect 27970 5705 31665 5725
rect 27480 5150 27520 5160
rect 27480 5130 27490 5150
rect 27510 5140 27520 5150
rect 27510 5130 27570 5140
rect 27480 5120 27570 5130
rect 27500 5080 27570 5100
<< viali >>
rect 27490 5130 27510 5150
<< metal1 >>
rect 27480 5310 27500 5385
rect 27480 5220 27625 5310
rect 27480 5160 27500 5220
rect 27480 5150 27520 5160
rect 27480 5130 27490 5150
rect 27510 5130 27520 5150
rect 27480 5120 27520 5130
rect 22920 3510 23630 4515
rect 23990 4510 26925 4515
rect 23990 3985 26830 4510
rect 26915 3985 26925 4510
rect 23990 3980 26925 3985
rect 27150 4510 31365 4515
rect 27150 3985 27160 4510
rect 27245 3985 31365 4510
rect 27150 3980 31365 3985
rect 30995 15 31365 3980
rect 30995 -520 34065 15
rect 33425 -1080 33525 -1075
rect 33425 -1260 33480 -1080
rect 33520 -1260 33525 -1080
rect 33425 -1265 33525 -1260
rect 33695 -1330 34065 -520
rect 33255 -1520 34065 -1330
<< via1 >>
rect 26830 3985 26915 4510
rect 27160 3985 27245 4510
rect 33480 -1260 33520 -1080
<< metal2 >>
rect 22650 5035 27010 5050
rect 22650 4725 26920 5035
rect 27000 4725 27010 5035
rect 22650 4710 27010 4725
rect 27150 5035 31365 5050
rect 27150 4725 27160 5035
rect 27240 4725 31365 5035
rect 27150 4710 31365 4725
rect 26820 4510 26925 4515
rect 26820 3985 26830 4510
rect 26915 3985 26925 4510
rect 26820 3980 26925 3985
rect 27150 4510 27255 4515
rect 27150 3985 27160 4510
rect 27245 3985 27255 4510
rect 27150 3980 27255 3985
rect 30995 15 31365 4710
rect 30995 -520 34065 15
rect 33695 -1075 34065 -520
rect 33475 -1080 34065 -1075
rect 33475 -1260 33480 -1080
rect 33520 -1260 34065 -1080
rect 33475 -1265 34065 -1260
<< via2 >>
rect 26920 4725 27000 5035
rect 27160 4725 27240 5035
rect 26830 3985 26915 4510
rect 27160 3985 27245 4510
<< metal3 >>
rect 27010 5045 27150 5050
rect 26910 5035 27250 5045
rect 26910 4725 26920 5035
rect 27000 4725 27160 5035
rect 27240 4725 27250 5035
rect 26910 4715 27250 4725
rect 27010 4710 27150 4715
rect 26820 4510 27255 4515
rect 26820 3985 26830 4510
rect 26915 3985 27160 4510
rect 27245 3985 27255 4510
rect 26820 3980 27255 3985
use adc  adc_0
timestamp 1620756519
transform 1 0 8045 0 1 -4180
box -7870 -175 25410 3310
use mux2  mux2_0
timestamp 1620437679
transform 1 0 27555 0 1 5200
box 0 -120 415 525
use bandgap_ping_pong  bandgap_ping_pong_0
timestamp 1620756519
transform 1 0 255 0 1 5525
box -255 -5525 30590 5560
<< end >>
