* NGSPICE file created from /home/madvlsi/Documents/MADVLSI-Final_Project/layout/inverter.ext - technology: sky130A

.subckt home/madvlsi/Documents/MADVLSI-Final_Project/layout/inverter A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=5e+06u as=1e+12p ps=5e+06u w=2e+06u l=150000u
.ends

