magic
tech sky130A
magscale 1 2
timestamp 1620691900
<< poly >>
rect -12860 6600 -12200 6630
rect -12860 5980 -12830 6600
rect -12230 6510 -12200 6600
rect -12230 6480 -6020 6510
rect -6050 6370 -6020 6480
rect -13750 5960 -13670 5980
rect -13750 5930 -13730 5960
rect -13880 5920 -13730 5930
rect -13690 5920 -13670 5960
rect -13880 5900 -13670 5920
rect -12910 5960 -12830 5980
rect -12910 5920 -12890 5960
rect -12850 5920 -12830 5960
rect -12910 5900 -12830 5920
rect -13880 5210 -13850 5900
rect -6120 4980 -6040 5000
rect -6120 4940 -6100 4980
rect -6060 4940 -6040 4980
rect -6120 4920 -6040 4940
rect -15990 3790 -15910 3810
rect -15990 3750 -15970 3790
rect -15930 3750 -15910 3790
rect -15990 3730 -15910 3750
<< polycont >>
rect -13730 5920 -13690 5960
rect -12890 5920 -12850 5960
rect -6100 4940 -6060 4980
rect -15970 3750 -15930 3790
<< locali >>
rect -11930 6480 -6080 6520
rect -11930 5980 -11890 6480
rect -13750 5960 -13670 5980
rect -13750 5920 -13730 5960
rect -13690 5950 -13670 5960
rect -13000 5960 -12700 5980
rect -13690 5920 -13640 5950
rect -13750 5910 -13640 5920
rect -13000 5920 -12890 5960
rect -12850 5920 -12700 5960
rect -13750 5900 -13650 5910
rect -13000 5900 -12700 5920
rect -12030 5900 -11890 5980
rect -15950 3810 -15910 5310
rect -6120 5000 -6080 6480
rect -6120 4980 -6040 5000
rect -6120 4940 -6100 4980
rect -6060 4940 -6040 4980
rect -6120 4920 -6040 4940
rect -15990 3790 -15910 3810
rect -15990 3750 -15970 3790
rect -15930 3750 -15910 3790
rect -15990 3730 -15910 3750
rect 270 1530 370 2100
rect -310 1460 16780 1530
rect 16730 160 16780 1460
rect 16730 150 17150 160
rect 16730 120 17160 150
use adc_digital  adc_digital_0
timestamp 1620691900
transform 1 0 0 0 1 3330
box 0 -3330 50820 3290
use comparator  comparator_0
timestamp 1620691900
transform 1 0 -5550 0 1 -3460
box -510 4630 5250 9940
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620691900
transform 1 0 -15410 0 1 -4650
box -510 4630 9129 11080
use switch  switch_0
timestamp 1620266915
transform 1 0 -12530 0 1 5300
box -180 40 500 1250
use switch  switch_1
timestamp 1620266915
transform 1 0 -13490 0 1 5300
box -180 40 500 1250
<< end >>
