magic
tech sky130A
timestamp 1620710927
<< poly >>
rect -60 2575 -15 2585
rect -60 2555 -50 2575
rect -30 2570 -15 2575
rect -30 2555 -20 2570
rect -60 2545 -20 2555
rect -375 1850 -15 1860
rect -375 1830 -365 1850
rect -345 1845 -15 1850
rect -345 1830 -335 1845
rect -375 1820 -335 1830
<< polycont >>
rect -50 2555 -30 2575
rect -365 1830 -345 1850
<< xpolycontact >>
rect -295 1250 -95 1275
<< locali >>
rect -1900 3155 2965 3175
rect -1900 1970 -1880 3155
rect -60 2575 -20 2585
rect -60 2555 -50 2575
rect -30 2555 -20 2575
rect -60 2545 -20 2555
rect -1900 1935 -1680 1970
rect -330 1915 -115 1935
rect -40 1915 -20 2545
rect -1045 1895 -20 1915
rect -2750 1735 -2530 1755
rect -1260 1740 -1220 1750
rect -1260 1735 -1250 1740
rect -2750 1720 -1250 1735
rect -1230 1735 -1220 1740
rect -1045 1735 -1025 1895
rect -375 1850 -335 1860
rect -375 1830 -365 1850
rect -345 1830 -335 1850
rect -375 1820 -335 1830
rect -1230 1720 -1025 1735
rect -2750 1715 -1025 1720
rect -1260 1710 -1220 1715
rect -3700 1485 -2895 1505
rect -3115 1430 -2895 1485
rect -2765 1485 -1025 1505
rect -2765 1465 -2545 1485
rect -1790 1280 -1570 1485
rect -1045 1365 -1025 1485
rect -355 1365 -335 1820
rect -1045 1345 -335 1365
rect 2945 540 2965 3155
<< viali >>
rect -3090 1760 -2890 1785
rect -1250 1720 -1230 1740
rect -295 1250 -95 1275
<< metal1 >>
rect -3100 1785 -2880 1790
rect -3100 1760 -3090 1785
rect -2890 1760 -2880 1785
rect -3100 1695 -2880 1760
rect -1260 1745 -1220 1750
rect -1260 1715 -1255 1745
rect -1225 1715 -1220 1745
rect -1260 1710 -1220 1715
rect -3100 1675 -1785 1695
rect -1805 1320 -1785 1675
rect -460 1400 -420 1405
rect -460 1370 -455 1400
rect -425 1370 -420 1400
rect -460 1320 -420 1370
rect -1805 1300 -85 1320
rect -305 1275 -85 1300
rect -305 1250 -295 1275
rect -95 1250 -85 1275
rect -305 1145 -85 1250
rect -305 1120 110 1145
<< via1 >>
rect -1255 1740 -1225 1745
rect -1255 1720 -1250 1740
rect -1250 1720 -1230 1740
rect -1230 1720 -1225 1740
rect -1255 1715 -1225 1720
rect -455 1370 -425 1400
<< metal2 >>
rect -1260 1745 -1220 1750
rect -1260 1715 -1255 1745
rect -1225 1715 -1220 1745
rect -1260 1710 -1220 1715
rect -460 1400 -420 1405
rect -460 1370 -455 1400
rect -425 1370 -420 1400
rect -460 1365 -420 1370
<< via2 >>
rect -1255 1715 -1225 1745
rect -455 1370 -425 1400
<< metal3 >>
rect -625 1895 -460 2430
rect -1265 1750 -1215 1755
rect -1265 1710 -1260 1750
rect -1220 1710 -1215 1750
rect -1265 1705 -1215 1710
rect -460 1400 -420 1405
rect -460 1370 -455 1400
rect -425 1370 -420 1400
rect -460 1365 -420 1370
<< via3 >>
rect -1260 1745 -1220 1750
rect -1260 1715 -1255 1745
rect -1255 1715 -1225 1745
rect -1225 1715 -1220 1745
rect -1260 1710 -1220 1715
<< metal4 >>
rect -775 1755 -675 2745
rect -1265 1750 -675 1755
rect -1265 1710 -1260 1750
rect -1220 1710 -675 1750
rect -1265 1705 -675 1710
rect -775 1670 -675 1705
use m3cap50f  m3cap50f_1
timestamp 1620687492
transform 1 0 -875 0 1 2445
box -115 -15 415 515
use m3cap50f  m3cap50f_0
timestamp 1620687492
transform 1 0 -875 0 1 1380
box -115 -15 415 515
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620692581
transform 1 0 235 0 1 -2345
box -255 2315 4445 5470
use p-res8x20k  p-res8x20k_1
timestamp 1620701388
transform 0 -1 -2875 1 0 1755
box 0 -915 590 795
use p-res8x20k  p-res8x20k_0
timestamp 1620701388
transform 0 1 -2770 -1 0 1465
box 0 -915 590 795
use p-res6x20k  p-res6x20k_1
timestamp 1620355847
transform 0 -1 -1025 1 0 2020
box -85 -915 320 790
use p-res6x20k  p-res6x20k_0
timestamp 1620355847
transform 0 1 -875 -1 0 1195
box -85 -915 320 790
<< end >>
