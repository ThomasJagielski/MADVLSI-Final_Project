magic
tech sky130A
timestamp 1620266915
<< nwell >>
rect -90 345 250 590
<< nmos >>
rect -40 75 -25 175
rect 35 75 50 275
rect 110 75 125 175
<< pmos >>
rect -40 470 -25 570
rect 35 370 50 570
rect 110 470 125 570
<< ndiff >>
rect -15 260 35 275
rect -15 175 0 260
rect -65 75 -40 175
rect -25 90 0 175
rect 20 90 35 260
rect -25 75 35 90
rect 50 260 100 275
rect 50 90 65 260
rect 85 175 100 260
rect 85 90 110 175
rect 50 75 110 90
rect 125 75 150 175
<< pdiff >>
rect -65 470 -40 570
rect -25 555 35 570
rect -25 470 0 555
rect -15 385 0 470
rect 20 385 35 555
rect -15 370 35 385
rect 50 555 110 570
rect 50 385 65 555
rect 85 470 110 555
rect 125 470 150 570
rect 85 385 100 470
rect 50 370 100 385
<< ndiffc >>
rect 0 90 20 260
rect 65 90 85 260
<< pdiffc >>
rect 0 385 20 555
rect 65 385 85 555
<< psubdiff >>
rect 180 160 230 175
rect 180 90 195 160
rect 215 90 230 160
rect 180 75 230 90
<< nsubdiff >>
rect 180 555 230 570
rect 180 485 195 555
rect 215 485 230 555
rect 180 470 230 485
<< psubdiffcont >>
rect 195 90 215 160
<< nsubdiffcont >>
rect 195 485 215 555
<< poly >>
rect -90 615 125 625
rect -90 595 -80 615
rect -60 610 125 615
rect -60 595 -25 610
rect -90 585 -25 595
rect -40 570 -25 585
rect 35 570 50 585
rect 110 570 125 610
rect -40 455 -25 470
rect 35 355 50 370
rect -40 340 50 355
rect -40 175 -25 340
rect 110 330 125 470
rect 70 315 125 330
rect 70 305 85 315
rect 35 290 85 305
rect 35 275 50 290
rect 110 175 125 290
rect -40 60 -25 75
rect 35 60 50 75
rect -90 50 -25 60
rect -90 30 -80 50
rect -60 35 -25 50
rect 110 35 125 75
rect -60 30 125 35
rect -90 20 125 30
<< polycont >>
rect -80 595 -60 615
rect -80 30 -60 50
<< locali >>
rect -90 615 -50 625
rect -90 595 -80 615
rect -60 595 -50 615
rect -90 585 -50 595
rect -10 555 30 565
rect -10 385 0 555
rect 20 385 30 555
rect -10 340 30 385
rect -90 300 30 340
rect -10 260 30 300
rect -10 90 0 260
rect 20 90 30 260
rect -10 80 30 90
rect 55 555 95 565
rect 55 385 65 555
rect 85 385 95 555
rect 185 555 225 565
rect 185 485 195 555
rect 215 485 225 555
rect 185 475 225 485
rect 55 340 95 385
rect 55 300 250 340
rect 55 260 95 300
rect 55 90 65 260
rect 85 90 95 260
rect 55 80 95 90
rect 185 160 225 170
rect 185 90 195 160
rect 215 90 225 160
rect 185 80 225 90
rect -90 50 -50 60
rect -90 30 -80 50
rect -60 30 -50 50
rect -90 20 -50 30
<< labels >>
rlabel locali -90 320 -90 320 7 A
rlabel locali 250 320 250 320 3 B
rlabel locali -90 40 -90 40 7 nCLK
rlabel locali -90 605 -90 605 7 CLK
<< end >>
