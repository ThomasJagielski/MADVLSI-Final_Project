magic
tech sky130A
timestamp 1620573865
<< nwell >>
rect 805 1270 1150 1295
rect 785 1080 1150 1270
rect 805 1055 1150 1080
rect 1010 395 1145 635
<< poly >>
rect 925 670 1130 680
rect 90 660 130 670
rect 90 640 100 660
rect 120 640 130 660
rect 90 630 130 640
rect 925 650 935 670
rect 955 665 1100 670
rect 955 650 965 665
rect 925 640 965 650
rect 1090 650 1100 665
rect 1120 650 1130 670
rect 1090 640 1130 650
rect 925 630 940 640
rect 985 25 1025 35
rect 985 5 995 25
rect 1015 10 1025 25
rect 1090 25 1130 35
rect 1090 10 1100 25
rect 1015 5 1100 10
rect 1120 5 1130 25
rect 985 -5 1130 5
<< polycont >>
rect 100 640 120 660
rect 935 650 955 670
rect 1100 650 1120 670
rect 995 5 1015 25
rect 1100 5 1120 25
<< locali >>
rect 760 1355 1150 1375
rect 760 1310 1070 1330
rect 805 765 945 785
rect 90 670 115 765
rect 735 700 900 720
rect 90 660 130 670
rect 90 640 100 660
rect 120 640 130 660
rect 90 630 130 640
rect 880 610 900 700
rect 925 680 945 765
rect 925 670 965 680
rect 925 650 935 670
rect 955 650 965 670
rect 925 640 965 650
rect 985 25 1025 35
rect 985 5 995 25
rect 1015 5 1025 25
rect 985 -5 1025 5
rect 1045 -30 1070 1310
rect 1090 765 1145 785
rect 1090 680 1110 765
rect 1090 670 1130 680
rect 1090 650 1100 670
rect 1120 650 1130 670
rect 1090 640 1130 650
rect 1090 25 1130 35
rect 1090 5 1100 25
rect 1120 15 1130 25
rect 1120 5 1145 15
rect 1090 -5 1145 5
rect 1010 -50 1070 -30
<< metal1 >>
rect 785 1190 1150 1270
rect 785 1160 840 1190
rect 870 1160 1150 1190
rect 785 1080 1150 1160
rect 805 935 1150 1015
rect 805 905 840 935
rect 870 905 1150 935
rect 805 825 1150 905
rect 510 695 590 710
rect 510 665 535 695
rect 565 665 590 695
rect 510 610 590 665
rect 1010 420 1145 610
rect 30 320 60 325
rect 30 295 40 320
rect 1010 165 1145 355
<< via1 >>
rect 840 1160 870 1190
rect 840 905 870 935
rect 535 665 565 695
rect 40 290 70 320
<< metal2 >>
rect 510 1190 925 1265
rect 510 1160 840 1190
rect 870 1160 925 1190
rect 510 1085 925 1160
rect 510 695 590 1085
rect 510 665 535 695
rect 565 665 590 695
rect 510 645 590 665
rect 790 935 925 1010
rect 790 905 840 935
rect 870 905 925 935
rect 790 350 925 905
rect 0 320 925 350
rect 0 290 40 320
rect 70 290 925 320
rect 0 265 925 290
use dff_upper  dff_upper_0
timestamp 1620491527
transform 1 0 -5 0 1 700
box 0 0 810 695
use dff_lower  dff_lower_0
timestamp 1620491637
transform 1 0 -35 0 1 130
box 30 -200 1045 505
<< labels >>
rlabel space -5 920 -5 920 7 GND
rlabel space -5 1175 -5 1175 7 VDD
rlabel space -5 775 -5 775 7 D
rlabel space -5 1320 -5 1320 7 CLK
rlabel space -5 1365 -5 1365 7 preset
rlabel locali 1145 775 1145 775 3 Q
rlabel space -5 5 -5 5 7 clear
<< end >>
