magic
tech sky130A
timestamp 1620778513
<< poly >>
rect -160 10875 210 10885
rect -160 10855 -150 10875
rect -130 10870 180 10875
rect -130 10855 -120 10870
rect -160 10845 -120 10855
rect 170 10855 180 10870
rect 200 10855 210 10875
rect 170 10845 210 10855
rect -115 8715 -70 8730
rect -115 8695 -105 8715
rect -80 8695 -70 8715
rect -115 8685 -70 8695
rect 33410 5715 33510 5725
rect 33410 5695 33420 5715
rect 33440 5710 33510 5715
rect 33440 5695 33450 5710
rect 33410 5685 33450 5695
<< polycont >>
rect -150 10855 -130 10875
rect 180 10855 200 10875
rect -105 8695 -80 8715
rect 33420 5695 33440 5715
<< locali >>
rect -140 18005 10010 18025
rect -140 10885 -120 18005
rect -160 10875 -120 10885
rect -160 10855 -150 10875
rect -130 10855 -120 10875
rect -160 10845 -120 10855
rect -100 17965 5045 17985
rect -100 8730 -80 17965
rect 5025 17920 5045 17965
rect -60 17255 15 17275
rect -60 10985 -40 17255
rect -60 10945 140 10985
rect 170 10875 210 10885
rect 170 10855 180 10875
rect 200 10855 210 10875
rect 170 10845 210 10855
rect -115 8715 -70 8730
rect -115 8695 -105 8715
rect -80 8695 -70 8715
rect -115 8685 -70 8695
rect 27555 5745 33495 5765
rect 27555 5705 27575 5745
rect 27970 5715 33450 5725
rect 27970 5705 33420 5715
rect 33410 5695 33420 5705
rect 33440 5695 33450 5715
rect 33410 5685 33450 5695
rect 27480 5120 27575 5140
rect 27480 5100 27500 5120
rect 32120 -2475 32160 -2420
rect 33475 -2475 33495 5745
rect 32120 -2495 33495 -2475
<< viali >>
rect -105 8695 -80 8715
rect 27915 5230 27935 5300
<< metal1 >>
rect 10350 11610 31365 11805
rect -115 8720 -70 8730
rect -115 8690 -110 8720
rect -75 8690 -70 8720
rect -115 8685 -70 8690
rect 27970 5655 28175 5665
rect 27970 5485 27985 5655
rect 28160 5485 28175 5655
rect 27970 5475 28175 5485
rect 27105 5310 27565 5410
rect 27105 5220 27625 5310
rect 30995 4515 31365 11610
rect 22920 3510 23630 4515
rect 23990 3980 31365 4515
rect 30995 15 31365 3980
rect 30995 -520 34065 15
rect 33425 -1080 33525 -1075
rect 33425 -1260 33480 -1080
rect 33520 -1260 33525 -1080
rect 33425 -1265 33525 -1260
rect 33695 -1330 34065 -520
rect 33255 -1520 34065 -1330
<< via1 >>
rect -110 8715 -75 8720
rect -110 8695 -105 8715
rect -105 8695 -80 8715
rect -80 8695 -75 8715
rect -110 8690 -75 8695
rect 27985 5485 28160 5655
rect 33480 -1260 33520 -1080
<< metal2 >>
rect 10265 11890 31365 12080
rect -115 8725 -70 8730
rect -115 8690 -110 8725
rect -75 8690 -70 8725
rect -115 8685 -70 8690
rect 27970 5655 28175 5665
rect 27970 5485 27985 5655
rect 28160 5485 28175 5655
rect 27970 5475 28175 5485
rect 28010 5050 28175 5475
rect 30995 5050 31365 11890
rect 22650 5035 27010 5050
rect 22650 4725 26920 5035
rect 27000 4725 27010 5035
rect 22650 4710 27010 4725
rect 27150 5035 31365 5050
rect 27150 4725 27160 5035
rect 27240 4725 31365 5035
rect 27150 4710 31365 4725
rect 30995 15 31365 4710
rect 30995 -520 34065 15
rect 33695 -1075 34065 -520
rect 33475 -1080 34065 -1075
rect 33475 -1260 33480 -1080
rect 33520 -1260 34065 -1080
rect 33475 -1265 34065 -1260
<< via2 >>
rect -110 8720 -75 8725
rect -110 8690 -75 8720
rect 26920 4725 27000 5035
rect 27160 4725 27240 5035
<< metal3 >>
rect -120 8725 5 8730
rect -120 8690 -110 8725
rect -75 8690 5 8725
rect -120 8680 5 8690
rect 27010 5045 27150 5050
rect 26910 5035 27250 5045
rect 26910 4725 26920 5035
rect 27000 4725 27160 5035
rect 27240 4725 27250 5035
rect 26910 4715 27250 4725
rect 27010 4710 27150 4715
use adc  adc_0
timestamp 1620778513
transform 1 0 8045 0 1 -4180
box -7870 -175 25410 3310
use bandgap  bandgap_0
timestamp 1620778513
transform 1 0 2160 0 1 14430
box -2180 -3165 12605 3600
use bandgap_ping_pong  bandgap_ping_pong_0
timestamp 1620778513
transform 1 0 255 0 1 5525
box -250 -5525 30590 5560
use mux2  mux2_0
timestamp 1620437679
transform 1 0 27555 0 1 5200
box 0 -120 415 525
<< labels >>
rlabel space 4105 3225 4105 3225 7 Vnn2
rlabel space 4085 8705 4085 8705 7 Vnn
rlabel space 4125 7965 4125 7965 7 Vpp
rlabel space 4145 2485 4145 2485 7 Vpp2
rlabel space 1390 8990 1390 8990 7 net9
rlabel space 1410 3510 1410 3510 7 net12
<< end >>
