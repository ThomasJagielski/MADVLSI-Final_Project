magic
tech sky130A
timestamp 1620615203
<< poly >>
rect 375 685 415 695
rect 375 665 385 685
rect 405 665 415 685
rect 375 655 415 665
rect 160 620 200 630
rect 160 600 170 620
rect 190 600 200 620
rect 160 590 200 600
rect 390 590 405 655
<< polycont >>
rect 385 665 405 685
rect 170 600 190 620
<< locali >>
rect 375 685 415 695
rect 375 675 385 685
rect 0 665 385 675
rect 405 675 415 685
rect 405 665 1015 675
rect 0 655 1015 665
rect 0 620 1015 630
rect 0 610 170 620
rect 160 600 170 610
rect 190 610 1015 620
rect 190 600 200 610
rect 160 590 200 600
rect 0 65 120 85
rect 225 40 245 90
rect 390 85 395 105
rect 715 65 865 85
rect 225 20 430 40
use nand2  nand2_2
timestamp 1620490283
transform 1 0 865 0 1 60
box -120 -60 150 535
use nand2  nand2_0
timestamp 1620490283
transform 1 0 120 0 1 60
box -120 -60 150 535
use and2  and2_0
timestamp 1620615203
transform 1 0 540 0 1 105
box -270 -105 205 490
<< end >>
