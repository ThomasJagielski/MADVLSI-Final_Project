magic
tech sky130A
timestamp 1620697439
<< nbase >>
rect 1230 -1770 1270 -1720
<< nmos >>
rect 2475 -615 2775 -555
rect 2475 -860 2775 -800
rect 2475 -980 2775 -920
rect 2475 -1100 2775 -1040
rect 2475 -1220 2775 -1160
rect 2475 -1340 2775 -1280
rect 2475 -1460 2775 -1400
rect 2475 -1580 2775 -1520
rect 2475 -1700 2775 -1640
rect 2475 -1940 2775 -1880
rect 2475 -2060 2775 -2000
rect 2475 -2180 2775 -2120
rect 2475 -2300 2775 -2240
rect 2475 -2420 2775 -2360
rect 2475 -2540 2775 -2480
rect 2475 -2660 2775 -2600
rect 2475 -2780 2775 -2720
rect 2475 -3025 2775 -2965
<< ndiff >>
rect 2475 -555 2775 -495
rect 2475 -685 2775 -615
rect 2475 -800 2775 -740
rect 2475 -920 2775 -860
rect 2475 -1040 2775 -980
rect 2475 -1160 2775 -1100
rect 2475 -1280 2775 -1220
rect 2475 -1400 2775 -1340
rect 2475 -1520 2775 -1460
rect 2475 -1640 2775 -1580
rect 2475 -1760 2775 -1700
rect 2475 -1880 2775 -1820
rect 2475 -2000 2775 -1940
rect 2475 -2120 2775 -2060
rect 2475 -2240 2775 -2180
rect 2475 -2360 2775 -2300
rect 2475 -2480 2775 -2420
rect 2475 -2600 2775 -2540
rect 2475 -2720 2775 -2660
rect 2475 -2845 2775 -2780
rect 2475 -2965 2775 -2900
rect 2475 -3085 2775 -3025
<< psubdiff >>
rect 2130 -505 2430 -495
rect 2130 -545 2145 -505
rect 2415 -545 2430 -505
rect 2130 -555 2430 -545
<< psubdiffcont >>
rect 2145 -545 2415 -505
<< poly >>
rect 2845 -510 2990 -500
rect 2845 -530 2855 -510
rect 2875 -520 2990 -510
rect 2875 -530 2885 -520
rect 2845 -540 2885 -530
rect 2445 -615 2475 -555
rect 2775 -615 2790 -555
rect 2445 -800 2460 -615
rect 2445 -860 2475 -800
rect 2775 -860 2790 -800
rect 2445 -920 2460 -860
rect 2445 -980 2475 -920
rect 2775 -980 2790 -920
rect 2445 -1040 2460 -980
rect 2445 -1100 2475 -1040
rect 2775 -1100 2790 -1040
rect 2445 -1160 2460 -1100
rect 2445 -1220 2475 -1160
rect 2775 -1220 2790 -1160
rect 2885 -1215 2925 -1205
rect 2445 -1280 2460 -1220
rect 2885 -1235 2895 -1215
rect 2915 -1225 2925 -1215
rect 2915 -1235 2995 -1225
rect 2885 -1245 2995 -1235
rect 2445 -1340 2475 -1280
rect 2775 -1340 2790 -1280
rect 2445 -1400 2460 -1340
rect 2445 -1460 2475 -1400
rect 2775 -1460 2790 -1400
rect 2445 -1520 2460 -1460
rect 2445 -1580 2475 -1520
rect 2775 -1580 2790 -1520
rect 2445 -1640 2460 -1580
rect 2445 -1700 2475 -1640
rect 2775 -1700 2790 -1640
rect 2445 -1880 2460 -1700
rect 2445 -1940 2475 -1880
rect 2775 -1940 2790 -1880
rect 2445 -2000 2460 -1940
rect 2445 -2060 2475 -2000
rect 2775 -2060 2790 -2000
rect 2445 -2120 2460 -2060
rect 2445 -2180 2475 -2120
rect 2775 -2180 2790 -2120
rect 2445 -2240 2460 -2180
rect 2445 -2300 2475 -2240
rect 2775 -2300 2790 -2240
rect 2445 -2360 2460 -2300
rect 2445 -2420 2475 -2360
rect 2775 -2420 2790 -2360
rect 2445 -2480 2460 -2420
rect 2445 -2540 2475 -2480
rect 2775 -2540 2790 -2480
rect 2445 -2600 2460 -2540
rect 2445 -2660 2475 -2600
rect 2775 -2660 2790 -2600
rect 2445 -2720 2460 -2660
rect 2445 -2780 2475 -2720
rect 2775 -2780 2790 -2720
rect 2445 -2965 2460 -2780
rect 2430 -3025 2475 -2965
rect 2775 -3025 2790 -2965
rect 2430 -3120 2445 -3025
rect 2430 -3130 2470 -3120
rect 2430 -3150 2440 -3130
rect 2460 -3150 2470 -3130
rect 2430 -3160 2470 -3150
<< polycont >>
rect 2855 -530 2875 -510
rect 2895 -1235 2915 -1215
rect 2440 -3150 2460 -3130
<< locali >>
rect 2135 -505 2425 -495
rect 2135 -545 2145 -505
rect 2415 -545 2425 -505
rect 2135 -555 2425 -545
rect 2480 -510 2770 -500
rect 2480 -540 2490 -510
rect 2760 -540 2770 -510
rect 2480 -550 2770 -540
rect 2845 -510 2885 -500
rect 2845 -530 2855 -510
rect 2875 -530 2885 -510
rect 2845 -540 2885 -530
rect 2480 -630 2770 -625
rect 2480 -670 2490 -630
rect 2760 -670 2770 -630
rect 2480 -675 2770 -670
rect 2435 -795 2770 -740
rect 2435 -975 2455 -795
rect 2480 -915 2815 -865
rect 1305 -985 2455 -975
rect 1305 -995 2770 -985
rect 1405 -1080 1460 -1030
rect 2435 -1035 2770 -995
rect 2435 -1225 2455 -1035
rect 2795 -1105 2815 -915
rect 2480 -1155 2815 -1105
rect 2435 -1275 2770 -1225
rect 2435 -1465 2455 -1275
rect 2795 -1345 2815 -1155
rect 2480 -1395 2815 -1345
rect 2435 -1515 2770 -1465
rect 2435 -1705 2455 -1515
rect 2795 -1585 2815 -1395
rect 2480 -1635 2815 -1585
rect 2845 -1655 2865 -540
rect 2795 -1675 2865 -1655
rect 2885 -1215 2925 -1205
rect 2885 -1235 2895 -1215
rect 2915 -1235 2925 -1215
rect 2885 -1245 2925 -1235
rect 2435 -1755 2770 -1705
rect 2435 -1875 2770 -1825
rect 2435 -2065 2455 -1875
rect 2795 -1945 2815 -1675
rect 2480 -1995 2815 -1945
rect 2435 -2115 2770 -2065
rect 2435 -2305 2455 -2115
rect 2795 -2185 2815 -1995
rect 2480 -2195 2815 -2185
rect 2480 -2225 2490 -2195
rect 2760 -2225 2815 -2195
rect 2480 -2235 2815 -2225
rect 2435 -2355 2770 -2305
rect 1010 -2545 1965 -2525
rect 1010 -2600 1230 -2545
rect 1945 -3030 1965 -2545
rect 2435 -2545 2455 -2355
rect 2795 -2425 2815 -2235
rect 2480 -2475 2815 -2425
rect 2435 -2595 2770 -2545
rect 2435 -2785 2455 -2595
rect 2795 -2665 2815 -2475
rect 2480 -2715 2815 -2665
rect 2435 -2795 2770 -2785
rect 2435 -2830 2485 -2795
rect 2755 -2830 2770 -2795
rect 2435 -2835 2770 -2830
rect 2480 -2840 2770 -2835
rect 2480 -2915 2770 -2905
rect 2480 -2950 2490 -2915
rect 2760 -2950 2770 -2915
rect 2480 -2960 2770 -2950
rect 2885 -3030 2910 -1245
rect 1945 -3080 2910 -3030
rect 2430 -3130 2470 -3120
rect 2430 -3150 2440 -3130
rect 2460 -3140 2470 -3130
rect 5920 -3140 5940 -2525
rect 2460 -3150 5940 -3140
rect 2430 -3160 5940 -3150
<< viali >>
rect 2145 -545 2415 -505
rect 2490 -540 2760 -510
rect 2490 -670 2760 -630
rect 1285 -995 1305 -975
rect 2490 -2225 2760 -2195
rect 2485 -2830 2755 -2795
rect 2490 -2950 2760 -2915
<< metal1 >>
rect 785 -510 2045 -490
rect 785 -705 810 -510
rect 2025 -625 2045 -510
rect 2135 -505 2830 -495
rect 2135 -545 2145 -505
rect 2415 -510 2830 -505
rect 2415 -540 2490 -510
rect 2760 -540 2830 -510
rect 2415 -545 2830 -540
rect 2135 -555 2830 -545
rect 2025 -630 2770 -625
rect 2025 -670 2490 -630
rect 2760 -670 2770 -630
rect 2025 -675 2770 -670
rect 1275 -975 1315 -965
rect 1275 -995 1285 -975
rect 1305 -995 1315 -975
rect 1275 -1215 1315 -995
rect 1230 -1725 1270 -1720
rect 1230 -1755 1235 -1725
rect 1265 -1755 1270 -1725
rect 1230 -1760 1270 -1755
rect 2480 -2195 2775 -2185
rect 2480 -2225 2490 -2195
rect 2760 -2225 2775 -2195
rect 2480 -2235 2775 -2225
rect 2480 -2795 2770 -2785
rect 2480 -2830 2485 -2795
rect 2755 -2830 2770 -2795
rect 2480 -2840 2770 -2830
rect 2480 -2915 2770 -2905
rect 2480 -2950 2490 -2915
rect 2760 -2950 2770 -2915
rect 2480 -2960 2770 -2950
<< via1 >>
rect 2145 -545 2415 -505
rect 2490 -540 2760 -510
rect 1235 -1755 1265 -1725
rect 2490 -2225 2760 -2195
rect 2485 -2830 2755 -2795
rect 2490 -2950 2760 -2915
<< metal2 >>
rect 2135 -505 2830 -495
rect 2135 -545 2145 -505
rect 2415 -510 2830 -505
rect 2415 -540 2490 -510
rect 2760 -540 2830 -510
rect 2415 -545 2830 -540
rect 2135 -555 2830 -545
rect 2810 -615 2830 -555
rect 2810 -645 3070 -615
rect 1230 -1725 1270 -1720
rect 1230 -1755 1235 -1725
rect 1265 -1755 1270 -1725
rect 1230 -1990 1270 -1755
rect 1230 -2010 2095 -1990
rect 2075 -2175 2095 -2010
rect 2075 -2195 2775 -2175
rect 2480 -2225 2490 -2195
rect 2760 -2225 2775 -2195
rect 2480 -2235 2775 -2225
rect 2480 -2795 2770 -2785
rect 2480 -2830 2485 -2795
rect 2755 -2830 2770 -2795
rect 2480 -2905 2770 -2830
rect 2480 -2915 2835 -2905
rect 2480 -2950 2490 -2915
rect 2760 -2950 2835 -2915
rect 2480 -2955 2835 -2950
rect 2480 -2960 2770 -2955
rect 2805 -3105 2835 -2955
rect 3185 -3105 3235 -2860
rect 2805 -3130 3235 -3105
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620692581
transform 1 0 3239 0 1 -5433
box -255 2315 4445 5470
use bandgap_pnp  bandgap_pnp_0
timestamp 1620689662
transform 1 0 1075 0 1 -915
box -2000 -2240 1155 898
<< end >>
