magic
tech sky130A
magscale 1 2
timestamp 1619188432
<< obsli1 >>
rect 1104 1445 45632 46257
<< obsm1 >>
rect 474 484 46078 46436
<< metal2 >>
rect 2778 48092 2834 48892
rect 6918 48092 6974 48892
rect 11518 48092 11574 48892
rect 15658 48092 15714 48892
rect 20258 48092 20314 48892
rect 24398 48092 24454 48892
rect 28998 48092 29054 48892
rect 33138 48092 33194 48892
rect 37738 48092 37794 48892
rect 41878 48092 41934 48892
rect 46018 48092 46074 48892
rect 478 0 534 800
rect 4618 0 4674 800
rect 8758 0 8814 800
rect 13358 0 13414 800
rect 17498 0 17554 800
rect 22098 0 22154 800
rect 26238 0 26294 800
rect 30838 0 30894 800
rect 34978 0 35034 800
rect 39578 0 39634 800
rect 43718 0 43774 800
<< obsm2 >>
rect 480 48036 2722 48092
rect 2890 48036 6862 48092
rect 7030 48036 11462 48092
rect 11630 48036 15602 48092
rect 15770 48036 20202 48092
rect 20370 48036 24342 48092
rect 24510 48036 28942 48092
rect 29110 48036 33082 48092
rect 33250 48036 37682 48092
rect 37850 48036 41822 48092
rect 41990 48036 45962 48092
rect 480 856 46072 48036
rect 590 478 4562 856
rect 4730 478 8702 856
rect 8870 478 13302 856
rect 13470 478 17442 856
rect 17610 478 22042 856
rect 22210 478 26182 856
rect 26350 478 30782 856
rect 30950 478 34922 856
rect 35090 478 39522 856
rect 39690 478 43662 856
rect 43830 478 46072 856
<< metal3 >>
rect 0 45568 800 45688
rect 45948 41488 46748 41608
rect 0 38768 800 38888
rect 45948 35368 46748 35488
rect 0 32648 800 32768
rect 45948 28568 46748 28688
rect 0 25848 800 25968
rect 45948 22448 46748 22568
rect 0 19728 800 19848
rect 45948 15648 46748 15768
rect 0 12928 800 13048
rect 45948 9528 46748 9648
rect 0 6808 800 6928
rect 45948 2728 46748 2848
<< obsm3 >>
rect 800 45768 45948 46273
rect 880 45488 45948 45768
rect 800 41688 45948 45488
rect 800 41408 45868 41688
rect 800 38968 45948 41408
rect 880 38688 45948 38968
rect 800 35568 45948 38688
rect 800 35288 45868 35568
rect 800 32848 45948 35288
rect 880 32568 45948 32848
rect 800 28768 45948 32568
rect 800 28488 45868 28768
rect 800 26048 45948 28488
rect 880 25768 45948 26048
rect 800 22648 45948 25768
rect 800 22368 45868 22648
rect 800 19928 45948 22368
rect 880 19648 45948 19928
rect 800 15848 45948 19648
rect 800 15568 45868 15848
rect 800 13128 45948 15568
rect 880 12848 45948 13128
rect 800 9728 45948 12848
rect 800 9448 45868 9728
rect 800 7008 45948 9448
rect 880 6728 45948 7008
rect 800 2928 45948 6728
rect 800 2648 45868 2928
rect 800 2143 45948 2648
<< metal4 >>
rect 4208 2128 4528 46288
rect 19568 2128 19888 46288
rect 34928 2128 35248 46288
<< obsm4 >>
rect 4659 4251 19488 44437
rect 19968 4251 34848 44437
rect 35328 4251 41341 44437
<< metal5 >>
rect 1104 35934 45632 36254
rect 1104 20616 45632 20936
rect 1104 5298 45632 5618
<< labels >>
rlabel metal3 s 0 6808 800 6928 6 DATA[0]
port 1 nsew signal output
rlabel metal2 s 20258 48092 20314 48892 6 DATA[10]
port 2 nsew signal output
rlabel metal2 s 28998 48092 29054 48892 6 DATA[11]
port 3 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 DATA[12]
port 4 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 DATA[13]
port 5 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 DATA[14]
port 6 nsew signal output
rlabel metal2 s 33138 48092 33194 48892 6 DATA[15]
port 7 nsew signal output
rlabel metal2 s 24398 48092 24454 48892 6 DATA[1]
port 8 nsew signal output
rlabel metal2 s 46018 48092 46074 48892 6 DATA[2]
port 9 nsew signal output
rlabel metal2 s 41878 48092 41934 48892 6 DATA[3]
port 10 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 DATA[4]
port 11 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 DATA[5]
port 12 nsew signal output
rlabel metal2 s 11518 48092 11574 48892 6 DATA[6]
port 13 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 DATA[7]
port 14 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 DATA[8]
port 15 nsew signal output
rlabel metal3 s 45948 28568 46748 28688 6 DATA[9]
port 16 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 data_en
port 17 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 dec_rate[0]
port 18 nsew signal input
rlabel metal3 s 45948 22448 46748 22568 6 dec_rate[10]
port 19 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 dec_rate[11]
port 20 nsew signal input
rlabel metal2 s 478 0 534 800 6 dec_rate[12]
port 21 nsew signal input
rlabel metal3 s 45948 2728 46748 2848 6 dec_rate[13]
port 22 nsew signal input
rlabel metal3 s 45948 35368 46748 35488 6 dec_rate[14]
port 23 nsew signal input
rlabel metal3 s 45948 9528 46748 9648 6 dec_rate[15]
port 24 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 dec_rate[1]
port 25 nsew signal input
rlabel metal2 s 2778 48092 2834 48892 6 dec_rate[2]
port 26 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 dec_rate[3]
port 27 nsew signal input
rlabel metal2 s 15658 48092 15714 48892 6 dec_rate[4]
port 28 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 dec_rate[5]
port 29 nsew signal input
rlabel metal2 s 37738 48092 37794 48892 6 dec_rate[6]
port 30 nsew signal input
rlabel metal3 s 45948 15648 46748 15768 6 dec_rate[7]
port 31 nsew signal input
rlabel metal2 s 6918 48092 6974 48892 6 dec_rate[8]
port 32 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 dec_rate[9]
port 33 nsew signal input
rlabel metal3 s 45948 41488 46748 41608 6 mclk1
port 34 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 mdata1
port 35 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 reset
port 36 nsew signal input
rlabel metal4 s 34928 2128 35248 46288 6 VPWR
port 37 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 46288 6 VPWR
port 38 nsew power bidirectional
rlabel metal5 s 1104 35934 45632 36254 6 VPWR
port 39 nsew power bidirectional
rlabel metal5 s 1104 5298 45632 5618 6 VPWR
port 40 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 46288 6 VGND
port 41 nsew ground bidirectional
rlabel metal5 s 1104 20616 45632 20936 6 VGND
port 42 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 46748 48892
string LEFview TRUE
string GDS_FILE /openLANE_flow/designs/decimation_filter/runs/23-04_14-21/results/magic/decimation_filter.gds
string GDS_END 7784476
string GDS_START 549836
<< end >>

