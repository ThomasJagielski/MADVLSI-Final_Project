magic
tech sky130A
timestamp 1620604183
<< nwell >>
rect -105 1370 -65 1375
rect 1355 1135 1390 1375
rect -200 690 5 715
rect -200 500 10 690
rect 1220 615 1395 715
rect 1220 505 1390 615
rect -200 475 5 500
rect 1220 475 1395 505
<< poly >>
rect 125 1540 2335 1555
rect -105 1505 -65 1515
rect -105 1485 -95 1505
rect -75 1485 -65 1505
rect -105 1475 -65 1485
rect -80 1410 -65 1475
rect -105 1400 -65 1410
rect -105 1380 -95 1400
rect -75 1380 -65 1400
rect -105 1370 -65 1380
rect 125 1370 140 1540
rect 1525 1505 1565 1515
rect 1525 1485 1535 1505
rect 1555 1485 1565 1505
rect 1525 1475 1565 1485
rect 1065 1465 1105 1475
rect 1065 1445 1075 1465
rect 1095 1445 1105 1465
rect 1065 1435 1105 1445
rect 1090 840 1105 1435
rect 1550 1410 1565 1475
rect 2320 1370 2335 1540
rect 1090 825 1220 840
rect 1205 750 1220 825
rect 1290 810 1330 820
rect 1290 795 1300 810
rect 1265 790 1300 795
rect 1320 790 1330 810
rect 1265 780 1330 790
rect 1205 735 1230 750
rect 1215 115 1230 735
rect 1265 155 1280 780
rect 1315 745 1355 755
rect 1315 725 1325 745
rect 1345 730 1355 745
rect 1345 725 1490 730
rect 1315 715 1490 725
rect 1265 140 1470 155
rect 1215 105 1430 115
rect 1215 100 1400 105
rect 1390 85 1400 100
rect 1420 85 1430 105
rect 1390 75 1430 85
rect 1455 50 1470 140
rect 1275 40 1470 50
rect 1275 20 1285 40
rect 1305 30 1470 40
rect 1305 20 1315 30
rect 1275 10 1315 20
rect 1510 -15 1525 185
rect 1820 0 1860 10
rect 1820 -15 1830 0
rect 1510 -20 1830 -15
rect 1850 -20 1860 0
rect 1510 -30 1860 -20
<< polycont >>
rect -95 1485 -75 1505
rect -95 1380 -75 1400
rect 1535 1485 1555 1505
rect 1075 1445 1095 1465
rect 1300 790 1320 810
rect 1325 725 1345 745
rect 1400 85 1420 105
rect 1285 20 1305 40
rect 1830 -20 1850 0
<< locali >>
rect -105 1505 1565 1515
rect -105 1485 -95 1505
rect -75 1495 1535 1505
rect -75 1485 -65 1495
rect -105 1475 -65 1485
rect 1525 1485 1535 1495
rect 1555 1485 1565 1505
rect 1525 1475 1565 1485
rect 1065 1465 1105 1475
rect -200 1435 5 1455
rect 1065 1445 1075 1465
rect 1095 1445 1105 1465
rect 1065 1435 1105 1445
rect 1350 1435 1405 1455
rect -200 1400 -65 1410
rect -200 1390 -95 1400
rect -105 1380 -95 1390
rect -75 1380 -65 1400
rect -105 1370 -65 1380
rect -40 1390 15 1410
rect -40 1350 -15 1390
rect 1220 845 1250 865
rect 1310 820 1330 850
rect 1290 810 1330 820
rect 1290 790 1300 810
rect 1320 790 1330 810
rect 1350 825 1370 1435
rect 1350 805 1395 825
rect 1290 780 1330 790
rect 1160 755 1180 765
rect 1160 745 1355 755
rect 1160 735 1325 745
rect 1315 725 1325 735
rect 1345 725 1355 745
rect 1315 715 1355 725
rect 1375 635 1395 805
rect 1350 615 1395 635
rect 1350 95 1370 615
rect -200 75 30 95
rect 1220 75 1370 95
rect 1390 105 1430 115
rect 1390 85 1400 105
rect 1420 85 1430 105
rect 1390 75 1430 85
rect -200 30 30 50
rect 1275 40 1315 50
rect 1275 20 1285 40
rect 1305 20 1315 40
rect 1275 5 1315 20
rect 1820 0 2610 10
rect 1820 -20 1830 0
rect 1850 -10 2610 0
rect 1850 -20 1860 -10
rect 1820 -30 1860 -20
<< metal1 >>
rect 1355 1160 1390 1350
rect 1355 905 1405 1095
rect -200 500 10 690
rect 1220 615 1395 690
rect 1220 500 1390 615
rect -200 245 5 435
rect 1220 245 1390 435
use dff  dff_0
timestamp 1620594849
transform 1 0 10 0 1 80
box -5 -70 1215 1395
use inverter  inverter_0
timestamp 1620435323
transform 1 0 -80 0 1 765
box -120 80 85 610
use inverter  inverter_1
timestamp 1620435323
transform 1 0 1270 0 1 765
box -120 80 85 610
use dff  dff_1
timestamp 1620594849
transform 1 0 1395 0 1 80
box -5 -70 1215 1395
<< labels >>
rlabel locali -200 1445 -200 1445 7 preset
rlabel locali -200 1400 -200 1400 7 CLK
rlabel locali 1295 5 1295 5 5 Qnout
rlabel locali 2610 0 2610 0 3 Qout
rlabel locali -200 85 -200 85 7 clear
<< end >>
