magic
tech sky130A
timestamp 1620703657
<< metal3 >>
rect 220 1545 3570 1645
rect 220 995 320 1545
rect 3470 995 3570 1545
rect 220 895 3570 995
rect 220 345 320 895
rect 3470 345 3570 895
rect 220 245 970 345
rect 1520 245 2270 345
rect 2820 245 3570 345
<< metal4 >>
rect 220 1545 3570 1645
rect 220 995 320 1545
rect 3470 995 3570 1545
rect 220 895 3570 995
rect 220 345 320 895
rect 3470 345 3570 895
rect 220 245 970 345
rect 1520 245 2270 345
rect 2820 245 3570 345
use m3cap50f  m3cap50f_7
timestamp 1620703657
transform 1 0 120 0 1 695
box -115 -15 415 515
use m3cap50f  m3cap50f_8
timestamp 1620703657
transform 1 0 770 0 1 695
box -115 -15 415 515
use m3cap50f  m3cap50f_3
timestamp 1620703657
transform 1 0 1420 0 1 695
box -115 -15 415 515
use m3cap50f  m3cap50f_14
timestamp 1620703657
transform -1 0 2370 0 1 695
box -115 -15 415 515
use m3cap50f  m3cap50f_9
timestamp 1620703657
transform -1 0 3020 0 1 695
box -115 -15 415 515
use m3cap50f  m3cap50f_6
timestamp 1620703657
transform 1 0 120 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_5
timestamp 1620703657
transform 1 0 770 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_4
timestamp 1620703657
transform 1 0 1420 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_13
timestamp 1620703657
transform -1 0 2370 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_12
timestamp 1620703657
transform -1 0 3020 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_0
timestamp 1620703657
transform 1 0 120 0 1 45
box -115 -15 415 515
use m3cap50f  m3cap50f_17
timestamp 1620703657
transform -1 0 3670 0 1 45
box -115 -15 415 515
use m3cap50f  m3cap50f_16
timestamp 1620703657
transform -1 0 3020 0 1 45
box -115 -15 415 515
use m3cap50f  m3cap50f_15
timestamp 1620703657
transform -1 0 2370 0 1 45
box -115 -15 415 515
use m3cap50f  m3cap50f_2
timestamp 1620703657
transform 1 0 1420 0 1 45
box -115 -15 415 515
use m3cap50f  m3cap50f_1
timestamp 1620703657
transform 1 0 770 0 1 45
box -115 -15 415 515
use m3cap50f  m3cap50f_10
timestamp 1620703657
transform -1 0 3670 0 1 695
box -115 -15 415 515
use m3cap50f  m3cap50f_11
timestamp 1620703657
transform -1 0 3670 0 1 1345
box -115 -15 415 515
<< end >>
