magic
tech sky130A
timestamp 1620661380
<< nwell >>
rect 1220 1125 1245 1365
rect 2460 1125 2480 1365
rect 3700 1125 3720 1365
rect 4940 1125 4960 1365
rect 6180 1125 6200 1365
rect 7420 1125 7440 1365
rect 8660 1125 8680 1365
rect 1220 465 1245 705
rect 2460 680 2480 705
rect 3700 680 3720 705
rect 2460 490 2485 680
rect 3695 490 3720 680
rect 2460 465 2480 490
rect 3700 465 3720 490
rect 4940 680 4960 705
rect 6180 680 6200 705
rect 4940 490 4965 680
rect 6180 490 6205 680
rect 4940 465 4960 490
rect 6180 465 6200 490
rect 7420 465 7440 705
rect 8660 680 8680 705
rect 8660 490 8685 680
rect 8660 465 8680 490
<< poly >>
rect 95 1495 135 1505
rect 95 1475 105 1495
rect 125 1475 135 1495
rect 95 1465 135 1475
rect 1335 1495 1375 1505
rect 1335 1475 1345 1495
rect 1365 1475 1375 1495
rect 1335 1465 1375 1475
rect 2575 1495 2615 1505
rect 2575 1475 2585 1495
rect 2605 1475 2615 1495
rect 2575 1465 2615 1475
rect 3815 1495 3855 1505
rect 3815 1475 3825 1495
rect 3845 1475 3855 1495
rect 3815 1465 3855 1475
rect 5055 1495 5095 1505
rect 5055 1475 5065 1495
rect 5085 1475 5095 1495
rect 5055 1465 5095 1475
rect 6295 1495 6335 1505
rect 6295 1475 6305 1495
rect 6325 1475 6335 1495
rect 6295 1465 6335 1475
rect 7535 1495 7575 1505
rect 7535 1475 7545 1495
rect 7565 1475 7575 1495
rect 7535 1465 7575 1475
rect 8775 1495 8815 1505
rect 8775 1475 8785 1495
rect 8805 1475 8815 1495
rect 8775 1465 8815 1475
rect 120 1360 135 1465
rect 1360 1360 1375 1465
rect 2600 1360 2615 1465
rect 3840 1355 3855 1465
rect 5080 1360 5095 1465
rect 6320 1360 6335 1465
rect 7560 1360 7575 1465
rect 8800 1360 8815 1465
rect 1070 0 1085 175
rect 2310 0 2325 175
rect 3550 0 3565 175
rect 4790 0 4805 175
rect 6030 0 6045 175
rect 7270 0 7285 175
rect 8510 0 8525 175
rect 9750 0 9765 175
rect 1045 -10 1085 0
rect 1045 -30 1055 -10
rect 1075 -30 1085 -10
rect 1045 -40 1085 -30
rect 2285 -10 2325 0
rect 2285 -30 2295 -10
rect 2315 -30 2325 -10
rect 2285 -40 2325 -30
rect 3525 -10 3565 0
rect 3525 -30 3535 -10
rect 3555 -30 3565 -10
rect 3525 -40 3565 -30
rect 4765 -10 4805 0
rect 4765 -30 4775 -10
rect 4795 -30 4805 -10
rect 4765 -40 4805 -30
rect 6005 -10 6045 0
rect 6005 -30 6015 -10
rect 6035 -30 6045 -10
rect 6005 -40 6045 -30
rect 7245 -10 7285 0
rect 7245 -30 7255 -10
rect 7275 -30 7285 -10
rect 7245 -40 7285 -30
rect 8485 -10 8525 0
rect 8485 -30 8495 -10
rect 8515 -30 8525 -10
rect 8485 -40 8525 -30
rect 9725 -10 9765 0
rect 9725 -30 9735 -10
rect 9755 -30 9765 -10
rect 9725 -40 9765 -30
<< polycont >>
rect 105 1475 125 1495
rect 1345 1475 1365 1495
rect 2585 1475 2605 1495
rect 3825 1475 3845 1495
rect 5065 1475 5085 1495
rect 6305 1475 6325 1495
rect 7545 1475 7565 1495
rect 8785 1475 8805 1495
rect 1055 -30 1075 -10
rect 2295 -30 2315 -10
rect 3535 -30 3555 -10
rect 4775 -30 4795 -10
rect 6015 -30 6035 -10
rect 7255 -30 7275 -10
rect 8495 -30 8515 -10
rect 9735 -30 9755 -10
<< locali >>
rect 95 1495 135 1505
rect 95 1475 105 1495
rect 125 1475 135 1495
rect 95 1465 135 1475
rect 1335 1495 1375 1505
rect 1335 1475 1345 1495
rect 1365 1475 1375 1495
rect 1335 1465 1375 1475
rect 2575 1495 2615 1505
rect 2575 1475 2585 1495
rect 2605 1475 2615 1495
rect 2575 1465 2615 1475
rect 3815 1495 3855 1505
rect 3815 1475 3825 1495
rect 3845 1475 3855 1495
rect 3815 1465 3855 1475
rect 5055 1495 5095 1505
rect 5055 1475 5065 1495
rect 5085 1475 5095 1495
rect 5055 1465 5095 1475
rect 6295 1495 6335 1505
rect 6295 1475 6305 1495
rect 6325 1475 6335 1495
rect 6295 1465 6335 1475
rect 7535 1495 7575 1505
rect 7535 1475 7545 1495
rect 7565 1475 7575 1495
rect 7535 1465 7575 1475
rect 8775 1495 8815 1505
rect 8775 1475 8785 1495
rect 8805 1475 8815 1495
rect 8775 1465 8815 1475
rect 0 1425 15 1445
rect 1215 1425 1250 1445
rect 2420 1425 2490 1445
rect 3690 1425 3730 1445
rect 4925 1425 4980 1445
rect 6170 1425 6220 1445
rect 7400 1425 7455 1445
rect 8650 1425 8700 1445
rect 0 1380 15 1400
rect 1215 1380 1250 1400
rect 2455 1380 2490 1400
rect 3690 1380 3725 1400
rect 4930 1380 4965 1400
rect 6170 1380 6205 1400
rect 7415 1380 7450 1400
rect 8655 1380 8690 1400
rect 0 65 15 85
rect 1215 65 1250 85
rect 2455 65 2485 85
rect 3700 65 3730 85
rect 4930 65 4975 85
rect 6180 65 6205 85
rect 7415 65 7450 85
rect 8655 65 8690 85
rect 1215 20 1250 40
rect 2455 20 2485 40
rect 3695 20 3725 40
rect 4930 20 4975 40
rect 6180 20 6205 40
rect 7415 20 7450 40
rect 8650 20 8685 40
rect 1045 -10 1085 0
rect 1045 -30 1055 -10
rect 1075 -30 1085 -10
rect 1045 -40 1085 -30
rect 2285 -10 2325 0
rect 2285 -30 2295 -10
rect 2315 -30 2325 -10
rect 2285 -40 2325 -30
rect 3525 -10 3565 0
rect 3525 -30 3535 -10
rect 3555 -30 3565 -10
rect 3525 -40 3565 -30
rect 4765 -10 4805 0
rect 4765 -30 4775 -10
rect 4795 -30 4805 -10
rect 4765 -40 4805 -30
rect 6005 -10 6045 0
rect 6005 -30 6015 -10
rect 6035 -30 6045 -10
rect 6005 -40 6045 -30
rect 7245 -10 7285 0
rect 7245 -30 7255 -10
rect 7275 -30 7285 -10
rect 7245 -40 7285 -30
rect 8485 -10 8525 0
rect 8485 -30 8495 -10
rect 8515 -30 8525 -10
rect 8485 -40 8525 -30
rect 9725 -10 9765 0
rect 9725 -30 9735 -10
rect 9755 -30 9765 -10
rect 9725 -40 9765 -30
<< metal1 >>
rect 0 1150 20 1340
rect 1220 1150 1240 1340
rect 2460 1150 2480 1340
rect 3700 1150 3720 1340
rect 4940 1150 4960 1340
rect 6180 1150 6200 1340
rect 7420 1150 7440 1340
rect 8660 1150 8680 1340
rect 0 895 15 1085
rect 1220 895 1240 1085
rect 2460 895 2480 1085
rect 3700 895 3720 1085
rect 4940 895 4960 1085
rect 6180 895 6200 1085
rect 7420 895 7440 1085
rect 8660 895 8680 1085
rect 1220 490 1240 680
rect 2460 490 2485 680
rect 3695 490 3720 680
rect 4940 490 4965 680
rect 6180 490 6205 680
rect 7420 490 7440 680
rect 8660 490 8685 680
rect 1220 235 1240 425
rect 2460 235 2485 425
rect 3700 235 3725 425
rect 4940 235 4965 425
rect 6175 235 6205 425
rect 7420 235 7440 425
rect 8660 235 8685 425
use dff  dff_7
timestamp 1620615203
transform 1 0 8685 0 1 70
box -5 -70 1215 1395
use dff  dff_6
timestamp 1620615203
transform 1 0 7445 0 1 70
box -5 -70 1215 1395
use dff  dff_5
timestamp 1620615203
transform 1 0 6205 0 1 70
box -5 -70 1215 1395
use dff  dff_4
timestamp 1620615203
transform 1 0 4965 0 1 70
box -5 -70 1215 1395
use dff  dff_3
timestamp 1620615203
transform 1 0 3725 0 1 70
box -5 -70 1215 1395
use dff  dff_2
timestamp 1620615203
transform 1 0 2485 0 1 70
box -5 -70 1215 1395
use dff  dff_1
timestamp 1620615203
transform 1 0 1245 0 1 70
box -5 -70 1215 1395
use dff  dff_0
timestamp 1620615203
transform 1 0 5 0 1 70
box -5 -70 1215 1395
<< labels >>
rlabel locali 115 1505 115 1505 1 Q0
rlabel locali 1355 1505 1355 1505 1 Q1
rlabel locali 2595 1505 2595 1505 1 Q2
rlabel locali 3835 1505 3835 1505 1 Q3
rlabel locali 5075 1505 5075 1505 1 Q4
rlabel locali 6315 1505 6315 1505 1 Q5
rlabel locali 7555 1505 7555 1505 1 Q6
rlabel locali 8795 1505 8795 1505 1 Q7
rlabel locali 1065 -40 1065 -40 5 Qout0
rlabel locali 2305 -40 2305 -40 5 Qout1
rlabel locali 3545 -40 3545 -40 5 Qout2
rlabel locali 4785 -40 4785 -40 5 Qout3
rlabel locali 6025 -40 6025 -40 5 Qout4
rlabel locali 7265 -40 7265 -40 5 Qout5
rlabel locali 8505 -40 8505 -40 5 Qout6
rlabel locali 9745 -40 9745 -40 5 Qout7
rlabel locali 0 1435 0 1435 7 preset
rlabel locali 0 1390 0 1390 7 CLK
rlabel metal1 0 1245 0 1245 7 VDD
rlabel metal1 0 990 0 990 7 GND
rlabel locali 0 75 0 75 7 clear
<< end >>
