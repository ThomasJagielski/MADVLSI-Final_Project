magic
tech sky130A
timestamp 1620688219
<< metal3 >>
rect 220 1545 3320 1645
rect 220 1045 320 1545
rect 3220 1045 3320 1545
rect 220 945 3320 1045
rect 220 445 320 945
rect 3220 445 3320 945
rect 220 345 920 445
rect 1420 345 2120 445
rect 2620 345 3320 445
<< metal4 >>
rect 220 1545 3320 1645
rect 220 1045 320 1545
rect 3220 1045 3320 1545
rect 220 945 3320 1045
rect 220 445 320 945
rect 3220 445 3320 945
rect 220 345 920 445
rect 1420 345 2120 445
rect 2620 345 3320 445
use m3cap50f  m3cap50f_0
timestamp 1620687492
transform 1 0 120 0 1 145
box -115 -15 415 515
use m3cap50f  m3cap50f_1
timestamp 1620687492
transform 1 0 720 0 1 145
box -115 -15 415 515
use m3cap50f  m3cap50f_2
timestamp 1620687492
transform 1 0 1320 0 1 145
box -115 -15 415 515
use m3cap50f  m3cap50f_15
timestamp 1620687492
transform -1 0 2220 0 1 145
box -115 -15 415 515
use m3cap50f  m3cap50f_16
timestamp 1620687492
transform -1 0 2820 0 1 145
box -115 -15 415 515
use m3cap50f  m3cap50f_7
timestamp 1620687492
transform 1 0 120 0 1 745
box -115 -15 415 515
use m3cap50f  m3cap50f_8
timestamp 1620687492
transform 1 0 720 0 1 745
box -115 -15 415 515
use m3cap50f  m3cap50f_3
timestamp 1620687492
transform 1 0 1320 0 1 745
box -115 -15 415 515
use m3cap50f  m3cap50f_14
timestamp 1620687492
transform -1 0 2220 0 1 745
box -115 -15 415 515
use m3cap50f  m3cap50f_9
timestamp 1620687492
transform -1 0 2820 0 1 745
box -115 -15 415 515
use m3cap50f  m3cap50f_6
timestamp 1620687492
transform 1 0 120 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_5
timestamp 1620687492
transform 1 0 720 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_4
timestamp 1620687492
transform 1 0 1320 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_13
timestamp 1620687492
transform -1 0 2220 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_12
timestamp 1620687492
transform -1 0 2820 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_17
timestamp 1620687492
transform -1 0 3420 0 1 145
box -115 -15 415 515
use m3cap50f  m3cap50f_11
timestamp 1620687492
transform -1 0 3420 0 1 1345
box -115 -15 415 515
use m3cap50f  m3cap50f_10
timestamp 1620687492
transform -1 0 3420 0 1 745
box -115 -15 415 515
<< end >>
