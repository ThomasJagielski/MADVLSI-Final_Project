magic
tech sky130A
timestamp 1620350317
<< nwell >>
rect -120 295 150 535
<< nmos >>
rect 25 60 40 260
rect 65 60 80 260
<< pmos >>
rect 0 315 15 515
rect 65 315 80 515
<< ndiff >>
rect -25 245 25 260
rect -25 175 -10 245
rect 10 175 25 245
rect -25 145 25 175
rect -25 75 -10 145
rect 10 75 25 145
rect -25 60 25 75
rect 40 60 65 260
rect 80 245 130 260
rect 80 175 95 245
rect 115 175 130 245
rect 80 145 130 175
rect 80 75 95 145
rect 115 75 130 145
rect 80 60 130 75
<< pdiff >>
rect -50 500 0 515
rect -50 430 -35 500
rect -15 430 0 500
rect -50 400 0 430
rect -50 330 -35 400
rect -15 330 0 400
rect -50 315 0 330
rect 15 500 65 515
rect 15 430 30 500
rect 50 430 65 500
rect 15 400 65 430
rect 15 330 30 400
rect 50 330 65 400
rect 15 315 65 330
rect 80 500 130 515
rect 80 430 95 500
rect 115 430 130 500
rect 80 400 130 430
rect 80 330 95 400
rect 115 330 130 400
rect 80 315 130 330
<< ndiffc >>
rect -10 175 10 245
rect -10 75 10 145
rect 95 175 115 245
rect 95 75 115 145
<< pdiffc >>
rect -35 430 -15 500
rect -35 330 -15 400
rect 30 430 50 500
rect 30 330 50 400
rect 95 430 115 500
rect 95 330 115 400
<< psubdiff >>
rect -75 245 -25 260
rect -75 175 -60 245
rect -40 175 -25 245
rect -75 145 -25 175
rect -75 75 -60 145
rect -40 75 -25 145
rect -75 60 -25 75
<< nsubdiff >>
rect -100 500 -50 515
rect -100 430 -85 500
rect -65 430 -50 500
rect -100 400 -50 430
rect -100 330 -85 400
rect -65 330 -50 400
rect -100 315 -50 330
<< psubdiffcont >>
rect -60 175 -40 245
rect -60 75 -40 145
<< nsubdiffcont >>
rect -85 430 -65 500
rect -85 330 -65 400
<< poly >>
rect 0 515 15 530
rect 65 515 80 530
rect 0 285 15 315
rect 0 270 40 285
rect 25 260 40 270
rect 65 260 80 315
rect 25 45 40 60
rect 0 35 40 45
rect 0 15 10 35
rect 30 15 40 35
rect 0 5 40 15
rect 65 -20 80 60
rect 40 -30 80 -20
rect 40 -50 50 -30
rect 70 -50 80 -30
rect 40 -60 80 -50
<< polycont >>
rect 10 15 30 35
rect 50 -50 70 -30
<< locali >>
rect -95 500 -5 510
rect -95 430 -85 500
rect -65 430 -35 500
rect -15 430 -5 500
rect -95 400 -5 430
rect -95 330 -85 400
rect -65 330 -35 400
rect -15 330 -5 400
rect -95 320 -5 330
rect 20 500 60 510
rect 20 430 30 500
rect 50 430 60 500
rect 20 400 60 430
rect 20 330 30 400
rect 50 330 60 400
rect 20 320 60 330
rect 85 500 125 510
rect 85 430 95 500
rect 115 430 125 500
rect 85 400 125 430
rect 85 330 95 400
rect 115 330 125 400
rect 85 320 125 330
rect 40 255 60 320
rect -70 245 20 255
rect -70 175 -60 245
rect -40 175 -10 245
rect 10 175 20 245
rect 40 245 125 255
rect 40 235 95 245
rect -70 145 20 175
rect -70 75 -60 145
rect -40 75 -10 145
rect 10 75 20 145
rect -70 65 20 75
rect 85 175 95 235
rect 115 175 125 245
rect 85 145 125 175
rect 85 75 95 145
rect 115 75 125 145
rect 85 65 125 75
rect 0 35 40 45
rect 0 15 10 35
rect 30 15 40 35
rect 105 25 125 65
rect 0 5 40 15
rect 40 -30 80 -20
rect 40 -50 50 -30
rect 70 -50 80 -30
rect 40 -60 80 -50
<< viali >>
rect -85 430 -65 500
rect -35 430 -15 500
rect -85 330 -65 400
rect -35 330 -15 400
rect 95 430 115 500
rect 95 330 115 400
rect -60 175 -40 245
rect -10 175 10 245
rect -60 75 -40 145
rect -10 75 10 145
<< metal1 >>
rect -120 500 150 510
rect -120 430 -85 500
rect -65 430 -35 500
rect -15 430 95 500
rect 115 430 150 500
rect -120 400 150 430
rect -120 330 -85 400
rect -65 330 -35 400
rect -15 330 95 400
rect 115 330 150 400
rect -120 320 150 330
rect -120 245 150 255
rect -120 175 -60 245
rect -40 175 -10 245
rect 10 175 150 245
rect -120 145 150 175
rect -120 75 -60 145
rect -40 75 -10 145
rect 10 75 150 145
rect -120 65 150 75
<< labels >>
rlabel metal1 -120 160 -120 160 7 VN
port 5 w
rlabel metal1 -120 415 -120 415 7 VP
port 4 w
rlabel locali 0 35 0 35 7 A
port 1 w
rlabel locali 40 -30 40 -30 7 B
port 2 w
rlabel locali 125 35 125 35 3 Y
port 3 e
<< end >>
