magic
tech sky130A
timestamp 1620621831
<< nwell >>
rect 6280 1695 6305 1935
rect 9115 1910 9140 1935
rect 11945 1910 11970 1935
rect 14775 1910 14795 1935
rect 17605 1910 17630 1935
rect 9115 1720 9145 1910
rect 11945 1720 11975 1910
rect 14775 1720 14800 1910
rect 17605 1720 17625 1910
rect 9115 1695 9140 1720
rect 11945 1695 11970 1720
rect 14775 1695 14795 1720
rect 17605 1695 17630 1720
rect 20435 1695 20455 1935
rect 23265 1695 23290 1935
rect 26095 1695 26120 1935
rect 6270 1035 6325 1275
rect 9110 1035 9250 1275
rect 11945 1035 11970 1275
rect 14775 1035 14795 1275
rect 17605 1250 17630 1275
rect 17600 1060 17630 1250
rect 17605 1035 17630 1060
rect 20435 1035 20455 1275
rect 23265 1250 23285 1275
rect 23265 1060 23290 1250
rect 23265 1035 23285 1060
rect 26095 1035 26115 1275
<< poly >>
rect 6355 1405 6410 1420
rect 6255 705 6295 715
rect 6255 685 6265 705
rect 6285 685 6295 705
rect 6255 675 6295 685
rect 6355 550 6370 1405
rect 6330 540 6370 550
rect 6330 520 6340 540
rect 6360 520 6370 540
rect 6255 485 6270 515
rect 6330 510 6370 520
rect 9135 665 9175 675
rect 9135 645 9145 665
rect 9165 645 9175 665
rect 9135 635 9175 645
rect 9135 485 9150 635
rect 9255 570 9270 1405
rect 9230 560 9270 570
rect 9230 540 9240 560
rect 9260 540 9270 560
rect 9230 530 9270 540
rect 11965 665 12005 675
rect 11965 645 11975 665
rect 11995 645 12005 665
rect 11965 635 12005 645
rect 11965 485 11980 635
rect 12085 570 12100 1405
rect 12060 560 12100 570
rect 12060 540 12070 560
rect 12090 540 12100 560
rect 12060 530 12100 540
rect 14795 665 14835 675
rect 14795 645 14805 665
rect 14825 645 14835 665
rect 14795 635 14835 645
rect 14795 485 14810 635
rect 14915 570 14930 1405
rect 14890 560 14930 570
rect 14890 540 14900 560
rect 14920 540 14930 560
rect 14890 530 14930 540
rect 17625 665 17665 675
rect 17625 645 17635 665
rect 17655 645 17665 665
rect 17625 635 17665 645
rect 17625 485 17640 635
rect 17745 570 17760 1405
rect 17720 560 17760 570
rect 17720 540 17730 560
rect 17750 540 17760 560
rect 17720 530 17760 540
rect 20455 665 20495 675
rect 20455 645 20465 665
rect 20485 645 20495 665
rect 20455 635 20495 645
rect 20455 485 20470 635
rect 20575 570 20590 1410
rect 20550 560 20590 570
rect 20550 540 20560 560
rect 20580 540 20590 560
rect 20550 530 20590 540
rect 23285 665 23325 675
rect 23285 645 23295 665
rect 23315 645 23325 665
rect 23285 635 23325 645
rect 23285 485 23300 635
rect 23405 570 23420 1405
rect 23380 560 23420 570
rect 23380 540 23390 560
rect 23410 540 23420 560
rect 23380 530 23420 540
rect 26115 665 26155 675
rect 26115 645 26125 665
rect 26145 645 26155 665
rect 26115 635 26155 645
rect 26115 485 26130 635
rect 26235 570 26250 1405
rect 26210 560 26250 570
rect 26210 540 26220 560
rect 26240 540 26250 560
rect 26210 530 26250 540
rect 6255 470 26130 485
<< polycont >>
rect 6265 685 6285 705
rect 6340 520 6360 540
rect 9145 645 9165 665
rect 9240 540 9260 560
rect 11975 645 11995 665
rect 12070 540 12090 560
rect 14805 645 14825 665
rect 14900 540 14920 560
rect 17635 645 17655 665
rect 17730 540 17750 560
rect 20465 645 20485 665
rect 20560 540 20580 560
rect 23295 645 23315 665
rect 23390 540 23410 560
rect 26125 645 26145 665
rect 26220 540 26240 560
<< locali >>
rect 6305 2095 26135 2115
rect 6305 2075 6325 2095
rect 4990 2055 6325 2075
rect 4990 2015 5010 2055
rect 6305 2015 6325 2055
rect 4825 1995 5010 2015
rect 9135 1995 9155 2095
rect 11965 1995 11985 2095
rect 14795 2015 14815 2095
rect 17625 2015 17645 2095
rect 20455 2015 20475 2095
rect 23285 2000 23305 2095
rect 26115 2015 26135 2095
rect 6255 705 6295 715
rect 6255 685 6265 705
rect 6285 695 6295 705
rect 6285 685 6325 695
rect 6255 675 6325 685
rect 6305 655 6325 675
rect 9135 665 9175 675
rect 9135 645 9145 665
rect 9165 645 9175 665
rect 9135 635 9175 645
rect 11965 665 12005 675
rect 11965 645 11975 665
rect 11995 645 12005 665
rect 11965 635 12005 645
rect 14795 665 14835 675
rect 14795 645 14805 665
rect 14825 645 14835 665
rect 14795 635 14835 645
rect 17625 665 17665 675
rect 17625 645 17635 665
rect 17655 645 17665 665
rect 17625 635 17665 645
rect 20455 665 20495 675
rect 20455 645 20465 665
rect 20485 645 20495 665
rect 20455 635 20495 645
rect 23285 665 23325 675
rect 23285 645 23295 665
rect 23315 645 23325 665
rect 23285 635 23325 645
rect 26115 665 26155 675
rect 26115 645 26125 665
rect 26145 645 26155 665
rect 26115 635 26155 645
rect 6330 540 6370 550
rect 6330 520 6340 540
rect 6360 520 6370 540
rect 6330 505 6370 520
rect 4960 485 6370 505
rect 7800 490 7820 570
rect 9230 560 9270 570
rect 9230 540 9240 560
rect 9260 540 9270 560
rect 9230 530 9270 540
rect 9230 490 9250 530
rect 7800 470 9250 490
rect 10630 490 10650 565
rect 12060 560 12100 570
rect 12060 540 12070 560
rect 12090 540 12100 560
rect 12060 530 12100 540
rect 12060 490 12080 530
rect 10630 470 12080 490
rect 13460 490 13480 565
rect 14890 560 14930 570
rect 14890 540 14900 560
rect 14920 540 14930 560
rect 14890 530 14930 540
rect 14890 490 14910 530
rect 13460 470 14910 490
rect 16290 490 16310 570
rect 17720 560 17760 570
rect 17720 540 17730 560
rect 17750 540 17760 560
rect 17720 530 17760 540
rect 17720 490 17740 530
rect 16290 470 17740 490
rect 19120 490 19140 565
rect 20550 560 20590 570
rect 20550 540 20560 560
rect 20580 540 20590 560
rect 20550 530 20590 540
rect 20550 490 20570 530
rect 19120 470 20570 490
rect 21950 490 21970 565
rect 23380 560 23420 570
rect 23380 540 23390 560
rect 23410 540 23420 560
rect 23380 530 23420 540
rect 23380 490 23400 530
rect 21950 470 23400 490
rect 24780 490 24800 565
rect 26210 560 26250 570
rect 26210 540 26220 560
rect 26240 540 26250 560
rect 26210 530 26250 540
rect 26210 490 26230 530
rect 24780 470 26230 490
<< metal1 >>
rect 6285 1720 6320 1910
rect 9115 1720 9145 1910
rect 11945 1720 11975 1910
rect 14775 1720 14800 1910
rect 17605 1720 17625 1910
rect 20435 1720 20455 1910
rect 23265 1720 23285 1910
rect 26095 1720 26120 1910
rect 6285 1465 6320 1655
rect 9115 1465 9145 1655
rect 11945 1465 11975 1655
rect 14775 1465 14805 1655
rect 17605 1465 17630 1655
rect 20435 1465 20455 1655
rect 23265 1465 23290 1655
rect 26095 1465 26120 1655
rect 6290 1060 6355 1250
rect 9115 1060 9145 1250
rect 11945 1060 11975 1250
rect 14775 1060 14805 1250
rect 17600 1060 17625 1250
rect 20435 1060 20455 1250
rect 23265 1060 23290 1250
rect 26095 1060 26115 1250
rect 6280 805 6345 995
rect 9110 805 9140 995
rect 11945 805 11975 995
rect 14775 805 14805 995
rect 17605 805 17630 995
rect 20435 805 20455 995
rect 23265 805 23290 995
rect 26095 805 26120 995
use counter_bn  counter_bn_7
timestamp 1620615203
transform 1 0 26315 0 1 560
box -200 -30 2610 1555
use counter_bn  counter_bn_6
timestamp 1620615203
transform 1 0 23485 0 1 560
box -200 -30 2610 1555
use counter_bn  counter_bn_5
timestamp 1620615203
transform 1 0 20655 0 1 560
box -200 -30 2610 1555
use counter_bn  counter_bn_4
timestamp 1620615203
transform 1 0 17825 0 1 560
box -200 -30 2610 1555
use counter_bn  counter_bn_3
timestamp 1620615203
transform 1 0 14995 0 1 560
box -200 -30 2610 1555
use counter_bn  counter_bn_2
timestamp 1620615203
transform 1 0 12165 0 1 560
box -200 -30 2610 1555
use counter_b0  counter_b0_0
timestamp 1620615203
transform 1 0 3605 0 1 570
box -90 -90 2685 1505
use counter_bn  counter_bn_0
timestamp 1620615203
transform 1 0 6505 0 1 560
box -200 -30 2610 1555
use counter_bn  counter_bn_1
timestamp 1620615203
transform 1 0 9335 0 1 560
box -200 -30 2610 1555
<< end >>
