magic
tech sky130A
timestamp 1620350971
use nand2  nand2_2
timestamp 1620350317
transform 1 0 895 0 1 -30
box -120 -60 150 535
use nand2  nand2_1
timestamp 1620350317
transform 1 0 625 0 1 -30
box -120 -60 150 535
use inverter  inverter_0
timestamp 1620350801
transform 1 0 150 0 1 -105
box -120 80 85 610
use nand2  nand2_0
timestamp 1620350317
transform 1 0 355 0 1 -30
box -120 -60 150 535
<< end >>
