**.subckt bandgap_thomas_test
XQ2 GND GND Vbep GND sky130_fd_pr__pnp_05v0
XQ4[7] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ4[6] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ4[5] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ4[4] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ4[3] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ4[2] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ4[1] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ4[0] GND GND Vben GND sky130_fd_pr__pnp_05v0
XQ1 GND GND net2 GND sky130_fd_pr__pnp_05v0
XQ3 GND __UNCONNECTED_PIN__0 net1 GND sky130_fd_pr__pnp_05v0
XQ4 GND __UNCONNECTED_PIN__1 __UNCONNECTED_PIN__2 GND sky130_fd_pr__pnp_05v0
XQ5 GND __UNCONNECTED_PIN__3 __UNCONNECTED_PIN__4 GND sky130_fd_pr__pnp_05v0
XQ6 GND __UNCONNECTED_PIN__5 __UNCONNECTED_PIN__6 GND sky130_fd_pr__pnp_05v0
XQ7 GND __UNCONNECTED_PIN__7 __UNCONNECTED_PIN__8 GND sky130_fd_pr__pnp_05v0
XQ8 GND __UNCONNECTED_PIN__9 __UNCONNECTED_PIN__10 GND sky130_fd_pr__pnp_05v0
XQ9 GND __UNCONNECTED_PIN__11 __UNCONNECTED_PIN__12 GND sky130_fd_pr__pnp_05v0
XQ10 GND __UNCONNECTED_PIN__13 __UNCONNECTED_PIN__14 GND sky130_fd_pr__pnp_05v0
XQ11 GND __UNCONNECTED_PIN__15 __UNCONNECTED_PIN__16 GND sky130_fd_pr__pnp_05v0
XQ12 GND __UNCONNECTED_PIN__17 __UNCONNECTED_PIN__18 GND sky130_fd_pr__pnp_05v0
XQ13 GND __UNCONNECTED_PIN__19 __UNCONNECTED_PIN__20 GND sky130_fd_pr__pnp_05v0
XQ14 GND __UNCONNECTED_PIN__21 __UNCONNECTED_PIN__22 GND sky130_fd_pr__pnp_05v0
XQ15 GND __UNCONNECTED_PIN__23 __UNCONNECTED_PIN__24 GND sky130_fd_pr__pnp_05v0
XQ16 GND __UNCONNECTED_PIN__25 __UNCONNECTED_PIN__26 GND sky130_fd_pr__pnp_05v0
XQ17 GND __UNCONNECTED_PIN__27 __UNCONNECTED_PIN__28 GND sky130_fd_pr__pnp_05v0
XQ18 GND __UNCONNECTED_PIN__29 __UNCONNECTED_PIN__30 GND sky130_fd_pr__pnp_05v0
XQ19 GND __UNCONNECTED_PIN__31 __UNCONNECTED_PIN__32 GND sky130_fd_pr__pnp_05v0
XQ20 GND __UNCONNECTED_PIN__33 __UNCONNECTED_PIN__34 GND sky130_fd_pr__pnp_05v0
XQ21 GND __UNCONNECTED_PIN__35 __UNCONNECTED_PIN__36 GND sky130_fd_pr__pnp_05v0
XQ22 GND __UNCONNECTED_PIN__37 __UNCONNECTED_PIN__38 GND sky130_fd_pr__pnp_05v0
**.ends
.GLOBAL GND
** flattened .save nodes
.end
