magic
tech sky130A
magscale 1 2
timestamp 1619963137
<< viali >>
rect 4261 15045 4295 15079
rect 4445 14841 4479 14875
rect 13277 11577 13311 11611
rect 13461 11577 13495 11611
rect 9668 11305 9702 11339
rect 9873 11237 9907 11271
rect 1961 11169 1995 11203
rect 1777 11033 1811 11067
rect 9505 10965 9539 10999
rect 9689 10965 9723 10999
rect 10333 10761 10367 10795
rect 10793 10693 10827 10727
rect 6837 10557 6871 10591
rect 8953 10557 8987 10591
rect 10793 10557 10827 10591
rect 11069 10557 11103 10591
rect 7082 10489 7116 10523
rect 9220 10489 9254 10523
rect 8217 10421 8251 10455
rect 10977 10421 11011 10455
rect 6653 10217 6687 10251
rect 8217 10217 8251 10251
rect 11437 10217 11471 10251
rect 7481 10149 7515 10183
rect 6193 10081 6227 10115
rect 6469 10081 6503 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 7619 10081 7653 10115
rect 8217 10081 8251 10115
rect 8401 10081 8435 10115
rect 10324 10081 10358 10115
rect 6285 10013 6319 10047
rect 7757 10013 7791 10047
rect 10057 10013 10091 10047
rect 7113 9877 7147 9911
rect 9413 9673 9447 9707
rect 10609 9673 10643 9707
rect 10057 9605 10091 9639
rect 6837 9469 6871 9503
rect 7104 9469 7138 9503
rect 9229 9469 9263 9503
rect 9413 9469 9447 9503
rect 9965 9469 9999 9503
rect 10428 9469 10462 9503
rect 8217 9333 8251 9367
rect 10425 9333 10459 9367
rect 8033 9129 8067 9163
rect 10149 9129 10183 9163
rect 8125 8993 8159 9027
rect 10241 8993 10275 9027
rect 8585 8585 8619 8619
rect 8769 8381 8803 8415
rect 10241 7293 10275 7327
rect 8953 7157 8987 7191
rect 9689 4777 9723 4811
rect 9505 4641 9539 4675
rect 10793 3621 10827 3655
rect 8125 3553 8159 3587
rect 9965 3553 9999 3587
rect 10149 3553 10183 3587
rect 10701 3553 10735 3587
rect 10885 3553 10919 3587
rect 10241 3485 10275 3519
rect 8217 3349 8251 3383
rect 9781 3349 9815 3383
rect 7941 3145 7975 3179
rect 11161 3145 11195 3179
rect 9321 3009 9355 3043
rect 9781 3009 9815 3043
rect 9054 2941 9088 2975
rect 10037 2941 10071 2975
rect 1961 2533 1995 2567
rect 8033 2533 8067 2567
rect 13277 2533 13311 2567
rect 1777 2329 1811 2363
rect 7849 2329 7883 2363
rect 13461 2329 13495 2363
<< metal1 >>
rect 1104 15258 14168 15280
rect 1104 15206 3159 15258
rect 3211 15206 3223 15258
rect 3275 15206 3287 15258
rect 3339 15206 3351 15258
rect 3403 15206 7514 15258
rect 7566 15206 7578 15258
rect 7630 15206 7642 15258
rect 7694 15206 7706 15258
rect 7758 15206 11868 15258
rect 11920 15206 11932 15258
rect 11984 15206 11996 15258
rect 12048 15206 12060 15258
rect 12112 15206 14168 15258
rect 1104 15184 14168 15206
rect 3694 15036 3700 15088
rect 3752 15076 3758 15088
rect 4249 15079 4307 15085
rect 4249 15076 4261 15079
rect 3752 15048 4261 15076
rect 3752 15036 3758 15048
rect 4249 15045 4261 15048
rect 4295 15045 4307 15079
rect 4249 15039 4307 15045
rect 4430 14872 4436 14884
rect 4391 14844 4436 14872
rect 4430 14832 4436 14844
rect 4488 14832 4494 14884
rect 1104 14714 14168 14736
rect 1104 14662 5336 14714
rect 5388 14662 5400 14714
rect 5452 14662 5464 14714
rect 5516 14662 5528 14714
rect 5580 14662 9691 14714
rect 9743 14662 9755 14714
rect 9807 14662 9819 14714
rect 9871 14662 9883 14714
rect 9935 14662 14168 14714
rect 1104 14640 14168 14662
rect 1104 14170 14168 14192
rect 1104 14118 3159 14170
rect 3211 14118 3223 14170
rect 3275 14118 3287 14170
rect 3339 14118 3351 14170
rect 3403 14118 7514 14170
rect 7566 14118 7578 14170
rect 7630 14118 7642 14170
rect 7694 14118 7706 14170
rect 7758 14118 11868 14170
rect 11920 14118 11932 14170
rect 11984 14118 11996 14170
rect 12048 14118 12060 14170
rect 12112 14118 14168 14170
rect 1104 14096 14168 14118
rect 1104 13626 14168 13648
rect 1104 13574 5336 13626
rect 5388 13574 5400 13626
rect 5452 13574 5464 13626
rect 5516 13574 5528 13626
rect 5580 13574 9691 13626
rect 9743 13574 9755 13626
rect 9807 13574 9819 13626
rect 9871 13574 9883 13626
rect 9935 13574 14168 13626
rect 1104 13552 14168 13574
rect 1104 13082 14168 13104
rect 1104 13030 3159 13082
rect 3211 13030 3223 13082
rect 3275 13030 3287 13082
rect 3339 13030 3351 13082
rect 3403 13030 7514 13082
rect 7566 13030 7578 13082
rect 7630 13030 7642 13082
rect 7694 13030 7706 13082
rect 7758 13030 11868 13082
rect 11920 13030 11932 13082
rect 11984 13030 11996 13082
rect 12048 13030 12060 13082
rect 12112 13030 14168 13082
rect 1104 13008 14168 13030
rect 1104 12538 14168 12560
rect 1104 12486 5336 12538
rect 5388 12486 5400 12538
rect 5452 12486 5464 12538
rect 5516 12486 5528 12538
rect 5580 12486 9691 12538
rect 9743 12486 9755 12538
rect 9807 12486 9819 12538
rect 9871 12486 9883 12538
rect 9935 12486 14168 12538
rect 1104 12464 14168 12486
rect 1104 11994 14168 12016
rect 1104 11942 3159 11994
rect 3211 11942 3223 11994
rect 3275 11942 3287 11994
rect 3339 11942 3351 11994
rect 3403 11942 7514 11994
rect 7566 11942 7578 11994
rect 7630 11942 7642 11994
rect 7694 11942 7706 11994
rect 7758 11942 11868 11994
rect 11920 11942 11932 11994
rect 11984 11942 11996 11994
rect 12048 11942 12060 11994
rect 12112 11942 14168 11994
rect 1104 11920 14168 11942
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 13265 11611 13323 11617
rect 13265 11608 13277 11611
rect 11020 11580 13277 11608
rect 11020 11568 11026 11580
rect 13265 11577 13277 11580
rect 13311 11577 13323 11611
rect 13446 11608 13452 11620
rect 13407 11580 13452 11608
rect 13265 11571 13323 11577
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 1104 11450 14168 11472
rect 1104 11398 5336 11450
rect 5388 11398 5400 11450
rect 5452 11398 5464 11450
rect 5516 11398 5528 11450
rect 5580 11398 9691 11450
rect 9743 11398 9755 11450
rect 9807 11398 9819 11450
rect 9871 11398 9883 11450
rect 9935 11398 14168 11450
rect 1104 11376 14168 11398
rect 9656 11339 9714 11345
rect 9656 11305 9668 11339
rect 9702 11336 9714 11339
rect 10042 11336 10048 11348
rect 9702 11308 10048 11336
rect 9702 11305 9714 11308
rect 9656 11299 9714 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 9861 11271 9919 11277
rect 9861 11237 9873 11271
rect 9907 11268 9919 11271
rect 10962 11268 10968 11280
rect 9907 11240 10968 11268
rect 9907 11237 9919 11240
rect 9861 11231 9919 11237
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 1995 11172 2774 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 1762 11064 1768 11076
rect 1723 11036 1768 11064
rect 1762 11024 1768 11036
rect 1820 11024 1826 11076
rect 2746 11064 2774 11172
rect 2746 11036 9720 11064
rect 9214 10956 9220 11008
rect 9272 10996 9278 11008
rect 9692 11005 9720 11036
rect 9493 10999 9551 11005
rect 9493 10996 9505 10999
rect 9272 10968 9505 10996
rect 9272 10956 9278 10968
rect 9493 10965 9505 10968
rect 9539 10965 9551 10999
rect 9493 10959 9551 10965
rect 9677 10999 9735 11005
rect 9677 10965 9689 10999
rect 9723 10996 9735 10999
rect 10318 10996 10324 11008
rect 9723 10968 10324 10996
rect 9723 10965 9735 10968
rect 9677 10959 9735 10965
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 1104 10906 14168 10928
rect 1104 10854 3159 10906
rect 3211 10854 3223 10906
rect 3275 10854 3287 10906
rect 3339 10854 3351 10906
rect 3403 10854 7514 10906
rect 7566 10854 7578 10906
rect 7630 10854 7642 10906
rect 7694 10854 7706 10906
rect 7758 10854 11868 10906
rect 11920 10854 11932 10906
rect 11984 10854 11996 10906
rect 12048 10854 12060 10906
rect 12112 10854 14168 10906
rect 1104 10832 14168 10854
rect 10318 10792 10324 10804
rect 10279 10764 10324 10792
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 10778 10724 10784 10736
rect 10739 10696 10784 10724
rect 10778 10684 10784 10696
rect 10836 10684 10842 10736
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 8938 10588 8944 10600
rect 8899 10560 8944 10588
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10376 10560 10793 10588
rect 10376 10548 10382 10560
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 6638 10480 6644 10532
rect 6696 10520 6702 10532
rect 7070 10523 7128 10529
rect 7070 10520 7082 10523
rect 6696 10492 7082 10520
rect 6696 10480 6702 10492
rect 7070 10489 7082 10492
rect 7116 10489 7128 10523
rect 7070 10483 7128 10489
rect 9208 10523 9266 10529
rect 9208 10489 9220 10523
rect 9254 10520 9266 10523
rect 9398 10520 9404 10532
rect 9254 10492 9404 10520
rect 9254 10489 9266 10492
rect 9208 10483 9266 10489
rect 9398 10480 9404 10492
rect 9456 10480 9462 10532
rect 10042 10480 10048 10532
rect 10100 10520 10106 10532
rect 11072 10520 11100 10551
rect 10100 10492 11100 10520
rect 10100 10480 10106 10492
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 10962 10452 10968 10464
rect 10923 10424 10968 10452
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 1104 10362 14168 10384
rect 1104 10310 5336 10362
rect 5388 10310 5400 10362
rect 5452 10310 5464 10362
rect 5516 10310 5528 10362
rect 5580 10310 9691 10362
rect 9743 10310 9755 10362
rect 9807 10310 9819 10362
rect 9871 10310 9883 10362
rect 9935 10310 14168 10362
rect 1104 10288 14168 10310
rect 6638 10248 6644 10260
rect 6599 10220 6644 10248
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7742 10248 7748 10260
rect 7156 10220 7748 10248
rect 7156 10208 7162 10220
rect 7742 10208 7748 10220
rect 7800 10248 7806 10260
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 7800 10220 8217 10248
rect 7800 10208 7806 10220
rect 8205 10217 8217 10220
rect 8251 10217 8263 10251
rect 8205 10211 8263 10217
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 11020 10220 11437 10248
rect 11020 10208 11026 10220
rect 11425 10217 11437 10220
rect 11471 10217 11483 10251
rect 11425 10211 11483 10217
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 7469 10183 7527 10189
rect 7469 10180 7481 10183
rect 7248 10152 7481 10180
rect 7248 10140 7254 10152
rect 7469 10149 7481 10152
rect 7515 10180 7527 10183
rect 7515 10152 8248 10180
rect 7515 10149 7527 10152
rect 7469 10143 7527 10149
rect 8220 10124 8248 10152
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 4488 10084 6193 10112
rect 4488 10072 4494 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 7098 10112 7104 10124
rect 6503 10084 7104 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 6196 9976 6224 10075
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 7282 10112 7288 10124
rect 7243 10084 7288 10112
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 7607 10115 7665 10121
rect 7607 10081 7619 10115
rect 7653 10112 7665 10115
rect 8018 10112 8024 10124
rect 7653 10084 8024 10112
rect 7653 10081 7665 10084
rect 7607 10075 7665 10081
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 7392 10044 7420 10075
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8202 10112 8208 10124
rect 8115 10084 8208 10112
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 9214 10112 9220 10124
rect 8435 10084 9220 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 7742 10044 7748 10056
rect 6319 10016 7420 10044
rect 7703 10016 7748 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 7190 9976 7196 9988
rect 6196 9948 7196 9976
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 7392 9976 7420 10016
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 8404 9976 8432 10075
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 10312 10115 10370 10121
rect 10312 10081 10324 10115
rect 10358 10112 10370 10115
rect 10594 10112 10600 10124
rect 10358 10084 10600 10112
rect 10358 10081 10370 10084
rect 10312 10075 10370 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 8628 10016 10057 10044
rect 8628 10004 8634 10016
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 7392 9948 8432 9976
rect 7098 9908 7104 9920
rect 7059 9880 7104 9908
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 1104 9818 14168 9840
rect 1104 9766 3159 9818
rect 3211 9766 3223 9818
rect 3275 9766 3287 9818
rect 3339 9766 3351 9818
rect 3403 9766 7514 9818
rect 7566 9766 7578 9818
rect 7630 9766 7642 9818
rect 7694 9766 7706 9818
rect 7758 9766 11868 9818
rect 11920 9766 11932 9818
rect 11984 9766 11996 9818
rect 12048 9766 12060 9818
rect 12112 9766 14168 9818
rect 1104 9744 14168 9766
rect 9398 9704 9404 9716
rect 9359 9676 9404 9704
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 10594 9704 10600 9716
rect 10555 9676 10600 9704
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 10042 9636 10048 9648
rect 10003 9608 10048 9636
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 10778 9568 10784 9580
rect 9416 9540 10784 9568
rect 6822 9500 6828 9512
rect 6735 9472 6828 9500
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7098 9509 7104 9512
rect 7092 9500 7104 9509
rect 7059 9472 7104 9500
rect 7092 9463 7104 9472
rect 7098 9460 7104 9463
rect 7156 9460 7162 9512
rect 9214 9500 9220 9512
rect 9175 9472 9220 9500
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9416 9509 9444 9540
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 10416 9503 10474 9509
rect 10416 9469 10428 9503
rect 10462 9469 10474 9503
rect 10416 9463 10474 9469
rect 6840 9432 6868 9460
rect 8570 9432 8576 9444
rect 6840 9404 8576 9432
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 9968 9432 9996 9463
rect 10428 9432 10456 9463
rect 10962 9432 10968 9444
rect 9968 9404 10968 9432
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 8076 9336 8217 9364
rect 8076 9324 8082 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10100 9336 10425 9364
rect 10100 9324 10106 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 1104 9274 14168 9296
rect 1104 9222 5336 9274
rect 5388 9222 5400 9274
rect 5452 9222 5464 9274
rect 5516 9222 5528 9274
rect 5580 9222 9691 9274
rect 9743 9222 9755 9274
rect 9807 9222 9819 9274
rect 9871 9222 9883 9274
rect 9935 9222 14168 9274
rect 1104 9200 14168 9222
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 8021 9163 8079 9169
rect 8021 9160 8033 9163
rect 7340 9132 8033 9160
rect 7340 9120 7346 9132
rect 8021 9129 8033 9132
rect 8067 9129 8079 9163
rect 8021 9123 8079 9129
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10137 9163 10195 9169
rect 10137 9160 10149 9163
rect 10100 9132 10149 9160
rect 10100 9120 10106 9132
rect 10137 9129 10149 9132
rect 10183 9129 10195 9163
rect 10137 9123 10195 9129
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 8076 8996 8125 9024
rect 8076 8984 8082 8996
rect 8113 8993 8125 8996
rect 8159 8993 8171 9027
rect 8113 8987 8171 8993
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 10100 8996 10241 9024
rect 10100 8984 10106 8996
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 1104 8730 14168 8752
rect 1104 8678 3159 8730
rect 3211 8678 3223 8730
rect 3275 8678 3287 8730
rect 3339 8678 3351 8730
rect 3403 8678 7514 8730
rect 7566 8678 7578 8730
rect 7630 8678 7642 8730
rect 7694 8678 7706 8730
rect 7758 8678 11868 8730
rect 11920 8678 11932 8730
rect 11984 8678 11996 8730
rect 12048 8678 12060 8730
rect 12112 8678 14168 8730
rect 1104 8656 14168 8678
rect 8570 8616 8576 8628
rect 8531 8588 8576 8616
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 8754 8412 8760 8424
rect 8715 8384 8760 8412
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 1104 8186 14168 8208
rect 1104 8134 5336 8186
rect 5388 8134 5400 8186
rect 5452 8134 5464 8186
rect 5516 8134 5528 8186
rect 5580 8134 9691 8186
rect 9743 8134 9755 8186
rect 9807 8134 9819 8186
rect 9871 8134 9883 8186
rect 9935 8134 14168 8186
rect 1104 8112 14168 8134
rect 1104 7642 14168 7664
rect 1104 7590 3159 7642
rect 3211 7590 3223 7642
rect 3275 7590 3287 7642
rect 3339 7590 3351 7642
rect 3403 7590 7514 7642
rect 7566 7590 7578 7642
rect 7630 7590 7642 7642
rect 7694 7590 7706 7642
rect 7758 7590 11868 7642
rect 11920 7590 11932 7642
rect 11984 7590 11996 7642
rect 12048 7590 12060 7642
rect 12112 7590 14168 7642
rect 1104 7568 14168 7590
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7324 10287 7327
rect 11054 7324 11060 7336
rect 10275 7296 11060 7324
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 8941 7191 8999 7197
rect 8941 7188 8953 7191
rect 8812 7160 8953 7188
rect 8812 7148 8818 7160
rect 8941 7157 8953 7160
rect 8987 7188 8999 7191
rect 9490 7188 9496 7200
rect 8987 7160 9496 7188
rect 8987 7157 8999 7160
rect 8941 7151 8999 7157
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 1104 7098 14168 7120
rect 1104 7046 5336 7098
rect 5388 7046 5400 7098
rect 5452 7046 5464 7098
rect 5516 7046 5528 7098
rect 5580 7046 9691 7098
rect 9743 7046 9755 7098
rect 9807 7046 9819 7098
rect 9871 7046 9883 7098
rect 9935 7046 14168 7098
rect 1104 7024 14168 7046
rect 1104 6554 14168 6576
rect 1104 6502 3159 6554
rect 3211 6502 3223 6554
rect 3275 6502 3287 6554
rect 3339 6502 3351 6554
rect 3403 6502 7514 6554
rect 7566 6502 7578 6554
rect 7630 6502 7642 6554
rect 7694 6502 7706 6554
rect 7758 6502 11868 6554
rect 11920 6502 11932 6554
rect 11984 6502 11996 6554
rect 12048 6502 12060 6554
rect 12112 6502 14168 6554
rect 1104 6480 14168 6502
rect 1104 6010 14168 6032
rect 1104 5958 5336 6010
rect 5388 5958 5400 6010
rect 5452 5958 5464 6010
rect 5516 5958 5528 6010
rect 5580 5958 9691 6010
rect 9743 5958 9755 6010
rect 9807 5958 9819 6010
rect 9871 5958 9883 6010
rect 9935 5958 14168 6010
rect 1104 5936 14168 5958
rect 1104 5466 14168 5488
rect 1104 5414 3159 5466
rect 3211 5414 3223 5466
rect 3275 5414 3287 5466
rect 3339 5414 3351 5466
rect 3403 5414 7514 5466
rect 7566 5414 7578 5466
rect 7630 5414 7642 5466
rect 7694 5414 7706 5466
rect 7758 5414 11868 5466
rect 11920 5414 11932 5466
rect 11984 5414 11996 5466
rect 12048 5414 12060 5466
rect 12112 5414 14168 5466
rect 1104 5392 14168 5414
rect 1104 4922 14168 4944
rect 1104 4870 5336 4922
rect 5388 4870 5400 4922
rect 5452 4870 5464 4922
rect 5516 4870 5528 4922
rect 5580 4870 9691 4922
rect 9743 4870 9755 4922
rect 9807 4870 9819 4922
rect 9871 4870 9883 4922
rect 9935 4870 14168 4922
rect 1104 4848 14168 4870
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9306 4808 9312 4820
rect 8996 4780 9312 4808
rect 8996 4768 9002 4780
rect 9306 4768 9312 4780
rect 9364 4808 9370 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 9364 4780 9689 4808
rect 9364 4768 9370 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 9677 4771 9735 4777
rect 9490 4672 9496 4684
rect 9451 4644 9496 4672
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 1104 4378 14168 4400
rect 1104 4326 3159 4378
rect 3211 4326 3223 4378
rect 3275 4326 3287 4378
rect 3339 4326 3351 4378
rect 3403 4326 7514 4378
rect 7566 4326 7578 4378
rect 7630 4326 7642 4378
rect 7694 4326 7706 4378
rect 7758 4326 11868 4378
rect 11920 4326 11932 4378
rect 11984 4326 11996 4378
rect 12048 4326 12060 4378
rect 12112 4326 14168 4378
rect 1104 4304 14168 4326
rect 1104 3834 14168 3856
rect 1104 3782 5336 3834
rect 5388 3782 5400 3834
rect 5452 3782 5464 3834
rect 5516 3782 5528 3834
rect 5580 3782 9691 3834
rect 9743 3782 9755 3834
rect 9807 3782 9819 3834
rect 9871 3782 9883 3834
rect 9935 3782 14168 3834
rect 1104 3760 14168 3782
rect 10781 3655 10839 3661
rect 10781 3652 10793 3655
rect 10060 3624 10793 3652
rect 10060 3596 10088 3624
rect 10781 3621 10793 3624
rect 10827 3621 10839 3655
rect 10781 3615 10839 3621
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3584 10011 3587
rect 10042 3584 10048 3596
rect 9999 3556 10048 3584
rect 9999 3553 10011 3556
rect 9953 3547 10011 3553
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8128 3516 8156 3547
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 10183 3556 10701 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10689 3553 10701 3556
rect 10735 3553 10747 3587
rect 10689 3547 10747 3553
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3553 10931 3587
rect 10873 3547 10931 3553
rect 10152 3516 10180 3547
rect 7984 3488 10180 3516
rect 10229 3519 10287 3525
rect 7984 3476 7990 3488
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10888 3516 10916 3547
rect 11146 3516 11152 3528
rect 10275 3488 11152 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 8202 3380 8208 3392
rect 8163 3352 8208 3380
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3380 9827 3383
rect 9858 3380 9864 3392
rect 9815 3352 9864 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 1104 3290 14168 3312
rect 1104 3238 3159 3290
rect 3211 3238 3223 3290
rect 3275 3238 3287 3290
rect 3339 3238 3351 3290
rect 3403 3238 7514 3290
rect 7566 3238 7578 3290
rect 7630 3238 7642 3290
rect 7694 3238 7706 3290
rect 7758 3238 11868 3290
rect 11920 3238 11932 3290
rect 11984 3238 11996 3290
rect 12048 3238 12060 3290
rect 12112 3238 14168 3290
rect 1104 3216 14168 3238
rect 7926 3176 7932 3188
rect 7887 3148 7932 3176
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 11146 3176 11152 3188
rect 11107 3148 11152 3176
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9306 3000 9312 3012
rect 9364 3040 9370 3052
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 9364 3012 9781 3040
rect 9364 3000 9370 3012
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 9042 2975 9100 2981
rect 9042 2972 9054 2975
rect 8260 2944 9054 2972
rect 8260 2932 8266 2944
rect 9042 2941 9054 2944
rect 9088 2941 9100 2975
rect 9042 2935 9100 2941
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 10025 2975 10083 2981
rect 10025 2972 10037 2975
rect 9916 2944 10037 2972
rect 9916 2932 9922 2944
rect 10025 2941 10037 2944
rect 10071 2941 10083 2975
rect 10025 2935 10083 2941
rect 1104 2746 14168 2768
rect 1104 2694 5336 2746
rect 5388 2694 5400 2746
rect 5452 2694 5464 2746
rect 5516 2694 5528 2746
rect 5580 2694 9691 2746
rect 9743 2694 9755 2746
rect 9807 2694 9819 2746
rect 9871 2694 9883 2746
rect 9935 2694 14168 2746
rect 1104 2672 14168 2694
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 7834 2564 7840 2576
rect 1995 2536 7840 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8018 2564 8024 2576
rect 7979 2536 8024 2564
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 13265 2567 13323 2573
rect 13265 2564 13277 2567
rect 11204 2536 13277 2564
rect 11204 2524 11210 2536
rect 13265 2533 13277 2536
rect 13311 2533 13323 2567
rect 13265 2527 13323 2533
rect 474 2320 480 2372
rect 532 2360 538 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 532 2332 1777 2360
rect 532 2320 538 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 7834 2360 7840 2372
rect 7795 2332 7840 2360
rect 1765 2323 1823 2329
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 13446 2360 13452 2372
rect 13407 2332 13452 2360
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 1104 2202 14168 2224
rect 1104 2150 3159 2202
rect 3211 2150 3223 2202
rect 3275 2150 3287 2202
rect 3339 2150 3351 2202
rect 3403 2150 7514 2202
rect 7566 2150 7578 2202
rect 7630 2150 7642 2202
rect 7694 2150 7706 2202
rect 7758 2150 11868 2202
rect 11920 2150 11932 2202
rect 11984 2150 11996 2202
rect 12048 2150 12060 2202
rect 12112 2150 14168 2202
rect 1104 2128 14168 2150
<< via1 >>
rect 3159 15206 3211 15258
rect 3223 15206 3275 15258
rect 3287 15206 3339 15258
rect 3351 15206 3403 15258
rect 7514 15206 7566 15258
rect 7578 15206 7630 15258
rect 7642 15206 7694 15258
rect 7706 15206 7758 15258
rect 11868 15206 11920 15258
rect 11932 15206 11984 15258
rect 11996 15206 12048 15258
rect 12060 15206 12112 15258
rect 3700 15036 3752 15088
rect 4436 14875 4488 14884
rect 4436 14841 4445 14875
rect 4445 14841 4479 14875
rect 4479 14841 4488 14875
rect 4436 14832 4488 14841
rect 5336 14662 5388 14714
rect 5400 14662 5452 14714
rect 5464 14662 5516 14714
rect 5528 14662 5580 14714
rect 9691 14662 9743 14714
rect 9755 14662 9807 14714
rect 9819 14662 9871 14714
rect 9883 14662 9935 14714
rect 3159 14118 3211 14170
rect 3223 14118 3275 14170
rect 3287 14118 3339 14170
rect 3351 14118 3403 14170
rect 7514 14118 7566 14170
rect 7578 14118 7630 14170
rect 7642 14118 7694 14170
rect 7706 14118 7758 14170
rect 11868 14118 11920 14170
rect 11932 14118 11984 14170
rect 11996 14118 12048 14170
rect 12060 14118 12112 14170
rect 5336 13574 5388 13626
rect 5400 13574 5452 13626
rect 5464 13574 5516 13626
rect 5528 13574 5580 13626
rect 9691 13574 9743 13626
rect 9755 13574 9807 13626
rect 9819 13574 9871 13626
rect 9883 13574 9935 13626
rect 3159 13030 3211 13082
rect 3223 13030 3275 13082
rect 3287 13030 3339 13082
rect 3351 13030 3403 13082
rect 7514 13030 7566 13082
rect 7578 13030 7630 13082
rect 7642 13030 7694 13082
rect 7706 13030 7758 13082
rect 11868 13030 11920 13082
rect 11932 13030 11984 13082
rect 11996 13030 12048 13082
rect 12060 13030 12112 13082
rect 5336 12486 5388 12538
rect 5400 12486 5452 12538
rect 5464 12486 5516 12538
rect 5528 12486 5580 12538
rect 9691 12486 9743 12538
rect 9755 12486 9807 12538
rect 9819 12486 9871 12538
rect 9883 12486 9935 12538
rect 3159 11942 3211 11994
rect 3223 11942 3275 11994
rect 3287 11942 3339 11994
rect 3351 11942 3403 11994
rect 7514 11942 7566 11994
rect 7578 11942 7630 11994
rect 7642 11942 7694 11994
rect 7706 11942 7758 11994
rect 11868 11942 11920 11994
rect 11932 11942 11984 11994
rect 11996 11942 12048 11994
rect 12060 11942 12112 11994
rect 10968 11568 11020 11620
rect 13452 11611 13504 11620
rect 13452 11577 13461 11611
rect 13461 11577 13495 11611
rect 13495 11577 13504 11611
rect 13452 11568 13504 11577
rect 5336 11398 5388 11450
rect 5400 11398 5452 11450
rect 5464 11398 5516 11450
rect 5528 11398 5580 11450
rect 9691 11398 9743 11450
rect 9755 11398 9807 11450
rect 9819 11398 9871 11450
rect 9883 11398 9935 11450
rect 10048 11296 10100 11348
rect 10968 11228 11020 11280
rect 1768 11067 1820 11076
rect 1768 11033 1777 11067
rect 1777 11033 1811 11067
rect 1811 11033 1820 11067
rect 1768 11024 1820 11033
rect 9220 10956 9272 11008
rect 10324 10956 10376 11008
rect 3159 10854 3211 10906
rect 3223 10854 3275 10906
rect 3287 10854 3339 10906
rect 3351 10854 3403 10906
rect 7514 10854 7566 10906
rect 7578 10854 7630 10906
rect 7642 10854 7694 10906
rect 7706 10854 7758 10906
rect 11868 10854 11920 10906
rect 11932 10854 11984 10906
rect 11996 10854 12048 10906
rect 12060 10854 12112 10906
rect 10324 10795 10376 10804
rect 10324 10761 10333 10795
rect 10333 10761 10367 10795
rect 10367 10761 10376 10795
rect 10324 10752 10376 10761
rect 10784 10727 10836 10736
rect 10784 10693 10793 10727
rect 10793 10693 10827 10727
rect 10827 10693 10836 10727
rect 10784 10684 10836 10693
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 10324 10548 10376 10600
rect 6644 10480 6696 10532
rect 9404 10480 9456 10532
rect 10048 10480 10100 10532
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 5336 10310 5388 10362
rect 5400 10310 5452 10362
rect 5464 10310 5516 10362
rect 5528 10310 5580 10362
rect 9691 10310 9743 10362
rect 9755 10310 9807 10362
rect 9819 10310 9871 10362
rect 9883 10310 9935 10362
rect 6644 10251 6696 10260
rect 6644 10217 6653 10251
rect 6653 10217 6687 10251
rect 6687 10217 6696 10251
rect 6644 10208 6696 10217
rect 7104 10208 7156 10260
rect 7748 10208 7800 10260
rect 10968 10208 11020 10260
rect 7196 10140 7248 10192
rect 4436 10072 4488 10124
rect 7104 10072 7156 10124
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 8024 10072 8076 10124
rect 8208 10115 8260 10124
rect 8208 10081 8217 10115
rect 8217 10081 8251 10115
rect 8251 10081 8260 10115
rect 8208 10072 8260 10081
rect 7748 10047 7800 10056
rect 7196 9936 7248 9988
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 9220 10072 9272 10124
rect 10600 10072 10652 10124
rect 8576 10004 8628 10056
rect 7104 9911 7156 9920
rect 7104 9877 7113 9911
rect 7113 9877 7147 9911
rect 7147 9877 7156 9911
rect 7104 9868 7156 9877
rect 3159 9766 3211 9818
rect 3223 9766 3275 9818
rect 3287 9766 3339 9818
rect 3351 9766 3403 9818
rect 7514 9766 7566 9818
rect 7578 9766 7630 9818
rect 7642 9766 7694 9818
rect 7706 9766 7758 9818
rect 11868 9766 11920 9818
rect 11932 9766 11984 9818
rect 11996 9766 12048 9818
rect 12060 9766 12112 9818
rect 9404 9707 9456 9716
rect 9404 9673 9413 9707
rect 9413 9673 9447 9707
rect 9447 9673 9456 9707
rect 9404 9664 9456 9673
rect 10600 9707 10652 9716
rect 10600 9673 10609 9707
rect 10609 9673 10643 9707
rect 10643 9673 10652 9707
rect 10600 9664 10652 9673
rect 10048 9639 10100 9648
rect 10048 9605 10057 9639
rect 10057 9605 10091 9639
rect 10091 9605 10100 9639
rect 10048 9596 10100 9605
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7104 9503 7156 9512
rect 7104 9469 7138 9503
rect 7138 9469 7156 9503
rect 7104 9460 7156 9469
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 10784 9528 10836 9580
rect 8576 9392 8628 9444
rect 10968 9392 11020 9444
rect 8024 9324 8076 9376
rect 10048 9324 10100 9376
rect 5336 9222 5388 9274
rect 5400 9222 5452 9274
rect 5464 9222 5516 9274
rect 5528 9222 5580 9274
rect 9691 9222 9743 9274
rect 9755 9222 9807 9274
rect 9819 9222 9871 9274
rect 9883 9222 9935 9274
rect 7288 9120 7340 9172
rect 10048 9120 10100 9172
rect 8024 8984 8076 9036
rect 10048 8984 10100 9036
rect 3159 8678 3211 8730
rect 3223 8678 3275 8730
rect 3287 8678 3339 8730
rect 3351 8678 3403 8730
rect 7514 8678 7566 8730
rect 7578 8678 7630 8730
rect 7642 8678 7694 8730
rect 7706 8678 7758 8730
rect 11868 8678 11920 8730
rect 11932 8678 11984 8730
rect 11996 8678 12048 8730
rect 12060 8678 12112 8730
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 5336 8134 5388 8186
rect 5400 8134 5452 8186
rect 5464 8134 5516 8186
rect 5528 8134 5580 8186
rect 9691 8134 9743 8186
rect 9755 8134 9807 8186
rect 9819 8134 9871 8186
rect 9883 8134 9935 8186
rect 3159 7590 3211 7642
rect 3223 7590 3275 7642
rect 3287 7590 3339 7642
rect 3351 7590 3403 7642
rect 7514 7590 7566 7642
rect 7578 7590 7630 7642
rect 7642 7590 7694 7642
rect 7706 7590 7758 7642
rect 11868 7590 11920 7642
rect 11932 7590 11984 7642
rect 11996 7590 12048 7642
rect 12060 7590 12112 7642
rect 11060 7284 11112 7336
rect 8760 7148 8812 7200
rect 9496 7148 9548 7200
rect 5336 7046 5388 7098
rect 5400 7046 5452 7098
rect 5464 7046 5516 7098
rect 5528 7046 5580 7098
rect 9691 7046 9743 7098
rect 9755 7046 9807 7098
rect 9819 7046 9871 7098
rect 9883 7046 9935 7098
rect 3159 6502 3211 6554
rect 3223 6502 3275 6554
rect 3287 6502 3339 6554
rect 3351 6502 3403 6554
rect 7514 6502 7566 6554
rect 7578 6502 7630 6554
rect 7642 6502 7694 6554
rect 7706 6502 7758 6554
rect 11868 6502 11920 6554
rect 11932 6502 11984 6554
rect 11996 6502 12048 6554
rect 12060 6502 12112 6554
rect 5336 5958 5388 6010
rect 5400 5958 5452 6010
rect 5464 5958 5516 6010
rect 5528 5958 5580 6010
rect 9691 5958 9743 6010
rect 9755 5958 9807 6010
rect 9819 5958 9871 6010
rect 9883 5958 9935 6010
rect 3159 5414 3211 5466
rect 3223 5414 3275 5466
rect 3287 5414 3339 5466
rect 3351 5414 3403 5466
rect 7514 5414 7566 5466
rect 7578 5414 7630 5466
rect 7642 5414 7694 5466
rect 7706 5414 7758 5466
rect 11868 5414 11920 5466
rect 11932 5414 11984 5466
rect 11996 5414 12048 5466
rect 12060 5414 12112 5466
rect 5336 4870 5388 4922
rect 5400 4870 5452 4922
rect 5464 4870 5516 4922
rect 5528 4870 5580 4922
rect 9691 4870 9743 4922
rect 9755 4870 9807 4922
rect 9819 4870 9871 4922
rect 9883 4870 9935 4922
rect 8944 4768 8996 4820
rect 9312 4768 9364 4820
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 3159 4326 3211 4378
rect 3223 4326 3275 4378
rect 3287 4326 3339 4378
rect 3351 4326 3403 4378
rect 7514 4326 7566 4378
rect 7578 4326 7630 4378
rect 7642 4326 7694 4378
rect 7706 4326 7758 4378
rect 11868 4326 11920 4378
rect 11932 4326 11984 4378
rect 11996 4326 12048 4378
rect 12060 4326 12112 4378
rect 5336 3782 5388 3834
rect 5400 3782 5452 3834
rect 5464 3782 5516 3834
rect 5528 3782 5580 3834
rect 9691 3782 9743 3834
rect 9755 3782 9807 3834
rect 9819 3782 9871 3834
rect 9883 3782 9935 3834
rect 7932 3476 7984 3528
rect 10048 3544 10100 3596
rect 11152 3476 11204 3528
rect 8208 3383 8260 3392
rect 8208 3349 8217 3383
rect 8217 3349 8251 3383
rect 8251 3349 8260 3383
rect 8208 3340 8260 3349
rect 9864 3340 9916 3392
rect 3159 3238 3211 3290
rect 3223 3238 3275 3290
rect 3287 3238 3339 3290
rect 3351 3238 3403 3290
rect 7514 3238 7566 3290
rect 7578 3238 7630 3290
rect 7642 3238 7694 3290
rect 7706 3238 7758 3290
rect 11868 3238 11920 3290
rect 11932 3238 11984 3290
rect 11996 3238 12048 3290
rect 12060 3238 12112 3290
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 11152 3179 11204 3188
rect 11152 3145 11161 3179
rect 11161 3145 11195 3179
rect 11195 3145 11204 3179
rect 11152 3136 11204 3145
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 8208 2932 8260 2984
rect 9864 2932 9916 2984
rect 5336 2694 5388 2746
rect 5400 2694 5452 2746
rect 5464 2694 5516 2746
rect 5528 2694 5580 2746
rect 9691 2694 9743 2746
rect 9755 2694 9807 2746
rect 9819 2694 9871 2746
rect 9883 2694 9935 2746
rect 7840 2524 7892 2576
rect 8024 2567 8076 2576
rect 8024 2533 8033 2567
rect 8033 2533 8067 2567
rect 8067 2533 8076 2567
rect 8024 2524 8076 2533
rect 11152 2524 11204 2576
rect 480 2320 532 2372
rect 7840 2363 7892 2372
rect 7840 2329 7849 2363
rect 7849 2329 7883 2363
rect 7883 2329 7892 2363
rect 7840 2320 7892 2329
rect 13452 2363 13504 2372
rect 13452 2329 13461 2363
rect 13461 2329 13495 2363
rect 13495 2329 13504 2363
rect 13452 2320 13504 2329
rect 3159 2150 3211 2202
rect 3223 2150 3275 2202
rect 3287 2150 3339 2202
rect 3351 2150 3403 2202
rect 7514 2150 7566 2202
rect 7578 2150 7630 2202
rect 7642 2150 7694 2202
rect 7706 2150 7758 2202
rect 11868 2150 11920 2202
rect 11932 2150 11984 2202
rect 11996 2150 12048 2202
rect 12060 2150 12112 2202
<< metal2 >>
rect 3698 16635 3754 17435
rect 11058 16635 11114 17435
rect 3133 15260 3429 15280
rect 3189 15258 3213 15260
rect 3269 15258 3293 15260
rect 3349 15258 3373 15260
rect 3211 15206 3213 15258
rect 3275 15206 3287 15258
rect 3349 15206 3351 15258
rect 3189 15204 3213 15206
rect 3269 15204 3293 15206
rect 3349 15204 3373 15206
rect 3133 15184 3429 15204
rect 3712 15094 3740 16635
rect 7488 15260 7784 15280
rect 7544 15258 7568 15260
rect 7624 15258 7648 15260
rect 7704 15258 7728 15260
rect 7566 15206 7568 15258
rect 7630 15206 7642 15258
rect 7704 15206 7706 15258
rect 7544 15204 7568 15206
rect 7624 15204 7648 15206
rect 7704 15204 7728 15206
rect 7488 15184 7784 15204
rect 3700 15088 3752 15094
rect 3700 15030 3752 15036
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 3133 14172 3429 14192
rect 3189 14170 3213 14172
rect 3269 14170 3293 14172
rect 3349 14170 3373 14172
rect 3211 14118 3213 14170
rect 3275 14118 3287 14170
rect 3349 14118 3351 14170
rect 3189 14116 3213 14118
rect 3269 14116 3293 14118
rect 3349 14116 3373 14118
rect 3133 14096 3429 14116
rect 3133 13084 3429 13104
rect 3189 13082 3213 13084
rect 3269 13082 3293 13084
rect 3349 13082 3373 13084
rect 3211 13030 3213 13082
rect 3275 13030 3287 13082
rect 3349 13030 3351 13082
rect 3189 13028 3213 13030
rect 3269 13028 3293 13030
rect 3349 13028 3373 13030
rect 3133 13008 3429 13028
rect 3133 11996 3429 12016
rect 3189 11994 3213 11996
rect 3269 11994 3293 11996
rect 3349 11994 3373 11996
rect 3211 11942 3213 11994
rect 3275 11942 3287 11994
rect 3349 11942 3351 11994
rect 3189 11940 3213 11942
rect 3269 11940 3293 11942
rect 3349 11940 3373 11942
rect 3133 11920 3429 11940
rect 1768 11076 1820 11082
rect 1768 11018 1820 11024
rect 1780 10985 1808 11018
rect 1766 10976 1822 10985
rect 1766 10911 1822 10920
rect 3133 10908 3429 10928
rect 3189 10906 3213 10908
rect 3269 10906 3293 10908
rect 3349 10906 3373 10908
rect 3211 10854 3213 10906
rect 3275 10854 3287 10906
rect 3349 10854 3351 10906
rect 3189 10852 3213 10854
rect 3269 10852 3293 10854
rect 3349 10852 3373 10854
rect 3133 10832 3429 10852
rect 4448 10130 4476 14826
rect 5310 14716 5606 14736
rect 5366 14714 5390 14716
rect 5446 14714 5470 14716
rect 5526 14714 5550 14716
rect 5388 14662 5390 14714
rect 5452 14662 5464 14714
rect 5526 14662 5528 14714
rect 5366 14660 5390 14662
rect 5446 14660 5470 14662
rect 5526 14660 5550 14662
rect 5310 14640 5606 14660
rect 9665 14716 9961 14736
rect 9721 14714 9745 14716
rect 9801 14714 9825 14716
rect 9881 14714 9905 14716
rect 9743 14662 9745 14714
rect 9807 14662 9819 14714
rect 9881 14662 9883 14714
rect 9721 14660 9745 14662
rect 9801 14660 9825 14662
rect 9881 14660 9905 14662
rect 9665 14640 9961 14660
rect 7488 14172 7784 14192
rect 7544 14170 7568 14172
rect 7624 14170 7648 14172
rect 7704 14170 7728 14172
rect 7566 14118 7568 14170
rect 7630 14118 7642 14170
rect 7704 14118 7706 14170
rect 7544 14116 7568 14118
rect 7624 14116 7648 14118
rect 7704 14116 7728 14118
rect 7488 14096 7784 14116
rect 5310 13628 5606 13648
rect 5366 13626 5390 13628
rect 5446 13626 5470 13628
rect 5526 13626 5550 13628
rect 5388 13574 5390 13626
rect 5452 13574 5464 13626
rect 5526 13574 5528 13626
rect 5366 13572 5390 13574
rect 5446 13572 5470 13574
rect 5526 13572 5550 13574
rect 5310 13552 5606 13572
rect 9665 13628 9961 13648
rect 9721 13626 9745 13628
rect 9801 13626 9825 13628
rect 9881 13626 9905 13628
rect 9743 13574 9745 13626
rect 9807 13574 9819 13626
rect 9881 13574 9883 13626
rect 9721 13572 9745 13574
rect 9801 13572 9825 13574
rect 9881 13572 9905 13574
rect 9665 13552 9961 13572
rect 7488 13084 7784 13104
rect 7544 13082 7568 13084
rect 7624 13082 7648 13084
rect 7704 13082 7728 13084
rect 7566 13030 7568 13082
rect 7630 13030 7642 13082
rect 7704 13030 7706 13082
rect 7544 13028 7568 13030
rect 7624 13028 7648 13030
rect 7704 13028 7728 13030
rect 7488 13008 7784 13028
rect 5310 12540 5606 12560
rect 5366 12538 5390 12540
rect 5446 12538 5470 12540
rect 5526 12538 5550 12540
rect 5388 12486 5390 12538
rect 5452 12486 5464 12538
rect 5526 12486 5528 12538
rect 5366 12484 5390 12486
rect 5446 12484 5470 12486
rect 5526 12484 5550 12486
rect 5310 12464 5606 12484
rect 9665 12540 9961 12560
rect 9721 12538 9745 12540
rect 9801 12538 9825 12540
rect 9881 12538 9905 12540
rect 9743 12486 9745 12538
rect 9807 12486 9819 12538
rect 9881 12486 9883 12538
rect 9721 12484 9745 12486
rect 9801 12484 9825 12486
rect 9881 12484 9905 12486
rect 9665 12464 9961 12484
rect 7488 11996 7784 12016
rect 7544 11994 7568 11996
rect 7624 11994 7648 11996
rect 7704 11994 7728 11996
rect 7566 11942 7568 11994
rect 7630 11942 7642 11994
rect 7704 11942 7706 11994
rect 7544 11940 7568 11942
rect 7624 11940 7648 11942
rect 7704 11940 7728 11942
rect 7488 11920 7784 11940
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 5310 11452 5606 11472
rect 5366 11450 5390 11452
rect 5446 11450 5470 11452
rect 5526 11450 5550 11452
rect 5388 11398 5390 11450
rect 5452 11398 5464 11450
rect 5526 11398 5528 11450
rect 5366 11396 5390 11398
rect 5446 11396 5470 11398
rect 5526 11396 5550 11398
rect 5310 11376 5606 11396
rect 9665 11452 9961 11472
rect 9721 11450 9745 11452
rect 9801 11450 9825 11452
rect 9881 11450 9905 11452
rect 9743 11398 9745 11450
rect 9807 11398 9819 11450
rect 9881 11398 9883 11450
rect 9721 11396 9745 11398
rect 9801 11396 9825 11398
rect 9881 11396 9905 11398
rect 9665 11376 9961 11396
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 7488 10908 7784 10928
rect 7544 10906 7568 10908
rect 7624 10906 7648 10908
rect 7704 10906 7728 10908
rect 7566 10854 7568 10906
rect 7630 10854 7642 10906
rect 7704 10854 7706 10906
rect 7544 10852 7568 10854
rect 7624 10852 7648 10854
rect 7704 10852 7728 10854
rect 7488 10832 7784 10852
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 5310 10364 5606 10384
rect 5366 10362 5390 10364
rect 5446 10362 5470 10364
rect 5526 10362 5550 10364
rect 5388 10310 5390 10362
rect 5452 10310 5464 10362
rect 5526 10310 5528 10362
rect 5366 10308 5390 10310
rect 5446 10308 5470 10310
rect 5526 10308 5550 10310
rect 5310 10288 5606 10308
rect 6656 10266 6684 10474
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 3133 9820 3429 9840
rect 3189 9818 3213 9820
rect 3269 9818 3293 9820
rect 3349 9818 3373 9820
rect 3211 9766 3213 9818
rect 3275 9766 3287 9818
rect 3349 9766 3351 9818
rect 3189 9764 3213 9766
rect 3269 9764 3293 9766
rect 3349 9764 3373 9766
rect 3133 9744 3429 9764
rect 6840 9518 6868 10542
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7116 10130 7144 10202
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7208 9994 7236 10134
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9518 7144 9862
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 5310 9276 5606 9296
rect 5366 9274 5390 9276
rect 5446 9274 5470 9276
rect 5526 9274 5550 9276
rect 5388 9222 5390 9274
rect 5452 9222 5464 9274
rect 5526 9222 5528 9274
rect 5366 9220 5390 9222
rect 5446 9220 5470 9222
rect 5526 9220 5550 9222
rect 5310 9200 5606 9220
rect 7300 9178 7328 10066
rect 7760 10062 7788 10202
rect 8220 10130 8248 10406
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7488 9820 7784 9840
rect 7544 9818 7568 9820
rect 7624 9818 7648 9820
rect 7704 9818 7728 9820
rect 7566 9766 7568 9818
rect 7630 9766 7642 9818
rect 7704 9766 7706 9818
rect 7544 9764 7568 9766
rect 7624 9764 7648 9766
rect 7704 9764 7728 9766
rect 7488 9744 7784 9764
rect 8036 9382 8064 10066
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9450 8616 9998
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 8036 9042 8064 9318
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 3133 8732 3429 8752
rect 3189 8730 3213 8732
rect 3269 8730 3293 8732
rect 3349 8730 3373 8732
rect 3211 8678 3213 8730
rect 3275 8678 3287 8730
rect 3349 8678 3351 8730
rect 3189 8676 3213 8678
rect 3269 8676 3293 8678
rect 3349 8676 3373 8678
rect 3133 8656 3429 8676
rect 7488 8732 7784 8752
rect 7544 8730 7568 8732
rect 7624 8730 7648 8732
rect 7704 8730 7728 8732
rect 7566 8678 7568 8730
rect 7630 8678 7642 8730
rect 7704 8678 7706 8730
rect 7544 8676 7568 8678
rect 7624 8676 7648 8678
rect 7704 8676 7728 8678
rect 7488 8656 7784 8676
rect 5310 8188 5606 8208
rect 5366 8186 5390 8188
rect 5446 8186 5470 8188
rect 5526 8186 5550 8188
rect 5388 8134 5390 8186
rect 5452 8134 5464 8186
rect 5526 8134 5528 8186
rect 5366 8132 5390 8134
rect 5446 8132 5470 8134
rect 5526 8132 5550 8134
rect 5310 8112 5606 8132
rect 3133 7644 3429 7664
rect 3189 7642 3213 7644
rect 3269 7642 3293 7644
rect 3349 7642 3373 7644
rect 3211 7590 3213 7642
rect 3275 7590 3287 7642
rect 3349 7590 3351 7642
rect 3189 7588 3213 7590
rect 3269 7588 3293 7590
rect 3349 7588 3373 7590
rect 3133 7568 3429 7588
rect 7488 7644 7784 7664
rect 7544 7642 7568 7644
rect 7624 7642 7648 7644
rect 7704 7642 7728 7644
rect 7566 7590 7568 7642
rect 7630 7590 7642 7642
rect 7704 7590 7706 7642
rect 7544 7588 7568 7590
rect 7624 7588 7648 7590
rect 7704 7588 7728 7590
rect 7488 7568 7784 7588
rect 5310 7100 5606 7120
rect 5366 7098 5390 7100
rect 5446 7098 5470 7100
rect 5526 7098 5550 7100
rect 5388 7046 5390 7098
rect 5452 7046 5464 7098
rect 5526 7046 5528 7098
rect 5366 7044 5390 7046
rect 5446 7044 5470 7046
rect 5526 7044 5550 7046
rect 5310 7024 5606 7044
rect 3133 6556 3429 6576
rect 3189 6554 3213 6556
rect 3269 6554 3293 6556
rect 3349 6554 3373 6556
rect 3211 6502 3213 6554
rect 3275 6502 3287 6554
rect 3349 6502 3351 6554
rect 3189 6500 3213 6502
rect 3269 6500 3293 6502
rect 3349 6500 3373 6502
rect 3133 6480 3429 6500
rect 7488 6556 7784 6576
rect 7544 6554 7568 6556
rect 7624 6554 7648 6556
rect 7704 6554 7728 6556
rect 7566 6502 7568 6554
rect 7630 6502 7642 6554
rect 7704 6502 7706 6554
rect 7544 6500 7568 6502
rect 7624 6500 7648 6502
rect 7704 6500 7728 6502
rect 7488 6480 7784 6500
rect 5310 6012 5606 6032
rect 5366 6010 5390 6012
rect 5446 6010 5470 6012
rect 5526 6010 5550 6012
rect 5388 5958 5390 6010
rect 5452 5958 5464 6010
rect 5526 5958 5528 6010
rect 5366 5956 5390 5958
rect 5446 5956 5470 5958
rect 5526 5956 5550 5958
rect 5310 5936 5606 5956
rect 3133 5468 3429 5488
rect 3189 5466 3213 5468
rect 3269 5466 3293 5468
rect 3349 5466 3373 5468
rect 3211 5414 3213 5466
rect 3275 5414 3287 5466
rect 3349 5414 3351 5466
rect 3189 5412 3213 5414
rect 3269 5412 3293 5414
rect 3349 5412 3373 5414
rect 3133 5392 3429 5412
rect 7488 5468 7784 5488
rect 7544 5466 7568 5468
rect 7624 5466 7648 5468
rect 7704 5466 7728 5468
rect 7566 5414 7568 5466
rect 7630 5414 7642 5466
rect 7704 5414 7706 5466
rect 7544 5412 7568 5414
rect 7624 5412 7648 5414
rect 7704 5412 7728 5414
rect 7488 5392 7784 5412
rect 5310 4924 5606 4944
rect 5366 4922 5390 4924
rect 5446 4922 5470 4924
rect 5526 4922 5550 4924
rect 5388 4870 5390 4922
rect 5452 4870 5464 4922
rect 5526 4870 5528 4922
rect 5366 4868 5390 4870
rect 5446 4868 5470 4870
rect 5526 4868 5550 4870
rect 5310 4848 5606 4868
rect 3133 4380 3429 4400
rect 3189 4378 3213 4380
rect 3269 4378 3293 4380
rect 3349 4378 3373 4380
rect 3211 4326 3213 4378
rect 3275 4326 3287 4378
rect 3349 4326 3351 4378
rect 3189 4324 3213 4326
rect 3269 4324 3293 4326
rect 3349 4324 3373 4326
rect 3133 4304 3429 4324
rect 7488 4380 7784 4400
rect 7544 4378 7568 4380
rect 7624 4378 7648 4380
rect 7704 4378 7728 4380
rect 7566 4326 7568 4378
rect 7630 4326 7642 4378
rect 7704 4326 7706 4378
rect 7544 4324 7568 4326
rect 7624 4324 7648 4326
rect 7704 4324 7728 4326
rect 7488 4304 7784 4324
rect 5310 3836 5606 3856
rect 5366 3834 5390 3836
rect 5446 3834 5470 3836
rect 5526 3834 5550 3836
rect 5388 3782 5390 3834
rect 5452 3782 5464 3834
rect 5526 3782 5528 3834
rect 5366 3780 5390 3782
rect 5446 3780 5470 3782
rect 5526 3780 5550 3782
rect 5310 3760 5606 3780
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 3133 3292 3429 3312
rect 3189 3290 3213 3292
rect 3269 3290 3293 3292
rect 3349 3290 3373 3292
rect 3211 3238 3213 3290
rect 3275 3238 3287 3290
rect 3349 3238 3351 3290
rect 3189 3236 3213 3238
rect 3269 3236 3293 3238
rect 3349 3236 3373 3238
rect 3133 3216 3429 3236
rect 7488 3292 7784 3312
rect 7544 3290 7568 3292
rect 7624 3290 7648 3292
rect 7704 3290 7728 3292
rect 7566 3238 7568 3290
rect 7630 3238 7642 3290
rect 7704 3238 7706 3290
rect 7544 3236 7568 3238
rect 7624 3236 7648 3238
rect 7704 3236 7728 3238
rect 7488 3216 7784 3236
rect 7944 3194 7972 3470
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7944 2774 7972 3130
rect 5310 2748 5606 2768
rect 5366 2746 5390 2748
rect 5446 2746 5470 2748
rect 5526 2746 5550 2748
rect 5388 2694 5390 2746
rect 5452 2694 5464 2746
rect 5526 2694 5528 2746
rect 5366 2692 5390 2694
rect 5446 2692 5470 2694
rect 5526 2692 5550 2694
rect 5310 2672 5606 2692
rect 7852 2746 7972 2774
rect 7852 2582 7880 2746
rect 8036 2582 8064 8978
rect 8588 8634 8616 9386
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8772 7206 8800 8366
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8956 4826 8984 10542
rect 9232 10130 9260 10950
rect 10060 10538 10088 11290
rect 10980 11286 11008 11562
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10810 10364 10950
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10336 10606 10364 10746
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9232 9518 9260 10066
rect 9416 9722 9444 10474
rect 9665 10364 9961 10384
rect 9721 10362 9745 10364
rect 9801 10362 9825 10364
rect 9881 10362 9905 10364
rect 9743 10310 9745 10362
rect 9807 10310 9819 10362
rect 9881 10310 9883 10362
rect 9721 10308 9745 10310
rect 9801 10308 9825 10310
rect 9881 10308 9905 10310
rect 9665 10288 9961 10308
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 10060 9654 10088 10474
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10612 9722 10640 10066
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 10060 9382 10088 9590
rect 10796 9586 10824 10678
rect 10980 10470 11008 11222
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10266 11008 10406
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10980 9450 11008 10202
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9665 9276 9961 9296
rect 9721 9274 9745 9276
rect 9801 9274 9825 9276
rect 9881 9274 9905 9276
rect 9743 9222 9745 9274
rect 9807 9222 9819 9274
rect 9881 9222 9883 9274
rect 9721 9220 9745 9222
rect 9801 9220 9825 9222
rect 9881 9220 9905 9222
rect 9665 9200 9961 9220
rect 10060 9178 10088 9318
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9665 8188 9961 8208
rect 9721 8186 9745 8188
rect 9801 8186 9825 8188
rect 9881 8186 9905 8188
rect 9743 8134 9745 8186
rect 9807 8134 9819 8186
rect 9881 8134 9883 8186
rect 9721 8132 9745 8134
rect 9801 8132 9825 8134
rect 9881 8132 9905 8134
rect 9665 8112 9961 8132
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8220 2990 8248 3334
rect 9324 3058 9352 4762
rect 9508 4690 9536 7142
rect 9665 7100 9961 7120
rect 9721 7098 9745 7100
rect 9801 7098 9825 7100
rect 9881 7098 9905 7100
rect 9743 7046 9745 7098
rect 9807 7046 9819 7098
rect 9881 7046 9883 7098
rect 9721 7044 9745 7046
rect 9801 7044 9825 7046
rect 9881 7044 9905 7046
rect 9665 7024 9961 7044
rect 9665 6012 9961 6032
rect 9721 6010 9745 6012
rect 9801 6010 9825 6012
rect 9881 6010 9905 6012
rect 9743 5958 9745 6010
rect 9807 5958 9819 6010
rect 9881 5958 9883 6010
rect 9721 5956 9745 5958
rect 9801 5956 9825 5958
rect 9881 5956 9905 5958
rect 9665 5936 9961 5956
rect 9665 4924 9961 4944
rect 9721 4922 9745 4924
rect 9801 4922 9825 4924
rect 9881 4922 9905 4924
rect 9743 4870 9745 4922
rect 9807 4870 9819 4922
rect 9881 4870 9883 4922
rect 9721 4868 9745 4870
rect 9801 4868 9825 4870
rect 9881 4868 9905 4870
rect 9665 4848 9961 4868
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9665 3836 9961 3856
rect 9721 3834 9745 3836
rect 9801 3834 9825 3836
rect 9881 3834 9905 3836
rect 9743 3782 9745 3834
rect 9807 3782 9819 3834
rect 9881 3782 9883 3834
rect 9721 3780 9745 3782
rect 9801 3780 9825 3782
rect 9881 3780 9905 3782
rect 9665 3760 9961 3780
rect 10060 3602 10088 8978
rect 11072 7342 11100 16635
rect 11842 15260 12138 15280
rect 11898 15258 11922 15260
rect 11978 15258 12002 15260
rect 12058 15258 12082 15260
rect 11920 15206 11922 15258
rect 11984 15206 11996 15258
rect 12058 15206 12060 15258
rect 11898 15204 11922 15206
rect 11978 15204 12002 15206
rect 12058 15204 12082 15206
rect 11842 15184 12138 15204
rect 11842 14172 12138 14192
rect 11898 14170 11922 14172
rect 11978 14170 12002 14172
rect 12058 14170 12082 14172
rect 11920 14118 11922 14170
rect 11984 14118 11996 14170
rect 12058 14118 12060 14170
rect 11898 14116 11922 14118
rect 11978 14116 12002 14118
rect 12058 14116 12082 14118
rect 11842 14096 12138 14116
rect 11842 13084 12138 13104
rect 11898 13082 11922 13084
rect 11978 13082 12002 13084
rect 12058 13082 12082 13084
rect 11920 13030 11922 13082
rect 11984 13030 11996 13082
rect 12058 13030 12060 13082
rect 11898 13028 11922 13030
rect 11978 13028 12002 13030
rect 12058 13028 12082 13030
rect 11842 13008 12138 13028
rect 11842 11996 12138 12016
rect 11898 11994 11922 11996
rect 11978 11994 12002 11996
rect 12058 11994 12082 11996
rect 11920 11942 11922 11994
rect 11984 11942 11996 11994
rect 12058 11942 12060 11994
rect 11898 11940 11922 11942
rect 11978 11940 12002 11942
rect 12058 11940 12082 11942
rect 11842 11920 12138 11940
rect 13450 11656 13506 11665
rect 13450 11591 13452 11600
rect 13504 11591 13506 11600
rect 13452 11562 13504 11568
rect 11842 10908 12138 10928
rect 11898 10906 11922 10908
rect 11978 10906 12002 10908
rect 12058 10906 12082 10908
rect 11920 10854 11922 10906
rect 11984 10854 11996 10906
rect 12058 10854 12060 10906
rect 11898 10852 11922 10854
rect 11978 10852 12002 10854
rect 12058 10852 12082 10854
rect 11842 10832 12138 10852
rect 11842 9820 12138 9840
rect 11898 9818 11922 9820
rect 11978 9818 12002 9820
rect 12058 9818 12082 9820
rect 11920 9766 11922 9818
rect 11984 9766 11996 9818
rect 12058 9766 12060 9818
rect 11898 9764 11922 9766
rect 11978 9764 12002 9766
rect 12058 9764 12082 9766
rect 11842 9744 12138 9764
rect 11842 8732 12138 8752
rect 11898 8730 11922 8732
rect 11978 8730 12002 8732
rect 12058 8730 12082 8732
rect 11920 8678 11922 8730
rect 11984 8678 11996 8730
rect 12058 8678 12060 8730
rect 11898 8676 11922 8678
rect 11978 8676 12002 8678
rect 12058 8676 12082 8678
rect 11842 8656 12138 8676
rect 11842 7644 12138 7664
rect 11898 7642 11922 7644
rect 11978 7642 12002 7644
rect 12058 7642 12082 7644
rect 11920 7590 11922 7642
rect 11984 7590 11996 7642
rect 12058 7590 12060 7642
rect 11898 7588 11922 7590
rect 11978 7588 12002 7590
rect 12058 7588 12082 7590
rect 11842 7568 12138 7588
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11842 6556 12138 6576
rect 11898 6554 11922 6556
rect 11978 6554 12002 6556
rect 12058 6554 12082 6556
rect 11920 6502 11922 6554
rect 11984 6502 11996 6554
rect 12058 6502 12060 6554
rect 11898 6500 11922 6502
rect 11978 6500 12002 6502
rect 12058 6500 12082 6502
rect 11842 6480 12138 6500
rect 11842 5468 12138 5488
rect 11898 5466 11922 5468
rect 11978 5466 12002 5468
rect 12058 5466 12082 5468
rect 11920 5414 11922 5466
rect 11984 5414 11996 5466
rect 12058 5414 12060 5466
rect 11898 5412 11922 5414
rect 11978 5412 12002 5414
rect 12058 5412 12082 5414
rect 11842 5392 12138 5412
rect 11842 4380 12138 4400
rect 11898 4378 11922 4380
rect 11978 4378 12002 4380
rect 12058 4378 12082 4380
rect 11920 4326 11922 4378
rect 11984 4326 11996 4378
rect 12058 4326 12060 4378
rect 11898 4324 11922 4326
rect 11978 4324 12002 4326
rect 12058 4324 12082 4326
rect 11842 4304 12138 4324
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9876 2990 9904 3334
rect 11164 3194 11192 3470
rect 11842 3292 12138 3312
rect 11898 3290 11922 3292
rect 11978 3290 12002 3292
rect 12058 3290 12082 3292
rect 11920 3238 11922 3290
rect 11984 3238 11996 3290
rect 12058 3238 12060 3290
rect 11898 3236 11922 3238
rect 11978 3236 12002 3238
rect 12058 3236 12082 3238
rect 11842 3216 12138 3236
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9665 2748 9961 2768
rect 9721 2746 9745 2748
rect 9801 2746 9825 2748
rect 9881 2746 9905 2748
rect 9743 2694 9745 2746
rect 9807 2694 9819 2746
rect 9881 2694 9883 2746
rect 9721 2692 9745 2694
rect 9801 2692 9825 2694
rect 9881 2692 9905 2694
rect 9665 2672 9961 2692
rect 11164 2582 11192 3130
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 480 2372 532 2378
rect 480 2314 532 2320
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 492 800 520 2314
rect 3133 2204 3429 2224
rect 3189 2202 3213 2204
rect 3269 2202 3293 2204
rect 3349 2202 3373 2204
rect 3211 2150 3213 2202
rect 3275 2150 3287 2202
rect 3349 2150 3351 2202
rect 3189 2148 3213 2150
rect 3269 2148 3293 2150
rect 3349 2148 3373 2150
rect 3133 2128 3429 2148
rect 7488 2204 7784 2224
rect 7544 2202 7568 2204
rect 7624 2202 7648 2204
rect 7704 2202 7728 2204
rect 7566 2150 7568 2202
rect 7630 2150 7642 2202
rect 7704 2150 7706 2202
rect 7544 2148 7568 2150
rect 7624 2148 7648 2150
rect 7704 2148 7728 2150
rect 7488 2128 7784 2148
rect 7852 800 7880 2314
rect 11842 2204 12138 2224
rect 11898 2202 11922 2204
rect 11978 2202 12002 2204
rect 12058 2202 12082 2204
rect 11920 2150 11922 2202
rect 11984 2150 11996 2202
rect 12058 2150 12060 2202
rect 11898 2148 11922 2150
rect 11978 2148 12002 2150
rect 12058 2148 12082 2150
rect 11842 2128 12138 2148
rect 478 0 534 800
rect 7838 0 7894 800
rect 13464 785 13492 2314
rect 13450 776 13506 785
rect 13450 711 13506 720
<< via2 >>
rect 3133 15258 3189 15260
rect 3213 15258 3269 15260
rect 3293 15258 3349 15260
rect 3373 15258 3429 15260
rect 3133 15206 3159 15258
rect 3159 15206 3189 15258
rect 3213 15206 3223 15258
rect 3223 15206 3269 15258
rect 3293 15206 3339 15258
rect 3339 15206 3349 15258
rect 3373 15206 3403 15258
rect 3403 15206 3429 15258
rect 3133 15204 3189 15206
rect 3213 15204 3269 15206
rect 3293 15204 3349 15206
rect 3373 15204 3429 15206
rect 7488 15258 7544 15260
rect 7568 15258 7624 15260
rect 7648 15258 7704 15260
rect 7728 15258 7784 15260
rect 7488 15206 7514 15258
rect 7514 15206 7544 15258
rect 7568 15206 7578 15258
rect 7578 15206 7624 15258
rect 7648 15206 7694 15258
rect 7694 15206 7704 15258
rect 7728 15206 7758 15258
rect 7758 15206 7784 15258
rect 7488 15204 7544 15206
rect 7568 15204 7624 15206
rect 7648 15204 7704 15206
rect 7728 15204 7784 15206
rect 3133 14170 3189 14172
rect 3213 14170 3269 14172
rect 3293 14170 3349 14172
rect 3373 14170 3429 14172
rect 3133 14118 3159 14170
rect 3159 14118 3189 14170
rect 3213 14118 3223 14170
rect 3223 14118 3269 14170
rect 3293 14118 3339 14170
rect 3339 14118 3349 14170
rect 3373 14118 3403 14170
rect 3403 14118 3429 14170
rect 3133 14116 3189 14118
rect 3213 14116 3269 14118
rect 3293 14116 3349 14118
rect 3373 14116 3429 14118
rect 3133 13082 3189 13084
rect 3213 13082 3269 13084
rect 3293 13082 3349 13084
rect 3373 13082 3429 13084
rect 3133 13030 3159 13082
rect 3159 13030 3189 13082
rect 3213 13030 3223 13082
rect 3223 13030 3269 13082
rect 3293 13030 3339 13082
rect 3339 13030 3349 13082
rect 3373 13030 3403 13082
rect 3403 13030 3429 13082
rect 3133 13028 3189 13030
rect 3213 13028 3269 13030
rect 3293 13028 3349 13030
rect 3373 13028 3429 13030
rect 3133 11994 3189 11996
rect 3213 11994 3269 11996
rect 3293 11994 3349 11996
rect 3373 11994 3429 11996
rect 3133 11942 3159 11994
rect 3159 11942 3189 11994
rect 3213 11942 3223 11994
rect 3223 11942 3269 11994
rect 3293 11942 3339 11994
rect 3339 11942 3349 11994
rect 3373 11942 3403 11994
rect 3403 11942 3429 11994
rect 3133 11940 3189 11942
rect 3213 11940 3269 11942
rect 3293 11940 3349 11942
rect 3373 11940 3429 11942
rect 1766 10920 1822 10976
rect 3133 10906 3189 10908
rect 3213 10906 3269 10908
rect 3293 10906 3349 10908
rect 3373 10906 3429 10908
rect 3133 10854 3159 10906
rect 3159 10854 3189 10906
rect 3213 10854 3223 10906
rect 3223 10854 3269 10906
rect 3293 10854 3339 10906
rect 3339 10854 3349 10906
rect 3373 10854 3403 10906
rect 3403 10854 3429 10906
rect 3133 10852 3189 10854
rect 3213 10852 3269 10854
rect 3293 10852 3349 10854
rect 3373 10852 3429 10854
rect 5310 14714 5366 14716
rect 5390 14714 5446 14716
rect 5470 14714 5526 14716
rect 5550 14714 5606 14716
rect 5310 14662 5336 14714
rect 5336 14662 5366 14714
rect 5390 14662 5400 14714
rect 5400 14662 5446 14714
rect 5470 14662 5516 14714
rect 5516 14662 5526 14714
rect 5550 14662 5580 14714
rect 5580 14662 5606 14714
rect 5310 14660 5366 14662
rect 5390 14660 5446 14662
rect 5470 14660 5526 14662
rect 5550 14660 5606 14662
rect 9665 14714 9721 14716
rect 9745 14714 9801 14716
rect 9825 14714 9881 14716
rect 9905 14714 9961 14716
rect 9665 14662 9691 14714
rect 9691 14662 9721 14714
rect 9745 14662 9755 14714
rect 9755 14662 9801 14714
rect 9825 14662 9871 14714
rect 9871 14662 9881 14714
rect 9905 14662 9935 14714
rect 9935 14662 9961 14714
rect 9665 14660 9721 14662
rect 9745 14660 9801 14662
rect 9825 14660 9881 14662
rect 9905 14660 9961 14662
rect 7488 14170 7544 14172
rect 7568 14170 7624 14172
rect 7648 14170 7704 14172
rect 7728 14170 7784 14172
rect 7488 14118 7514 14170
rect 7514 14118 7544 14170
rect 7568 14118 7578 14170
rect 7578 14118 7624 14170
rect 7648 14118 7694 14170
rect 7694 14118 7704 14170
rect 7728 14118 7758 14170
rect 7758 14118 7784 14170
rect 7488 14116 7544 14118
rect 7568 14116 7624 14118
rect 7648 14116 7704 14118
rect 7728 14116 7784 14118
rect 5310 13626 5366 13628
rect 5390 13626 5446 13628
rect 5470 13626 5526 13628
rect 5550 13626 5606 13628
rect 5310 13574 5336 13626
rect 5336 13574 5366 13626
rect 5390 13574 5400 13626
rect 5400 13574 5446 13626
rect 5470 13574 5516 13626
rect 5516 13574 5526 13626
rect 5550 13574 5580 13626
rect 5580 13574 5606 13626
rect 5310 13572 5366 13574
rect 5390 13572 5446 13574
rect 5470 13572 5526 13574
rect 5550 13572 5606 13574
rect 9665 13626 9721 13628
rect 9745 13626 9801 13628
rect 9825 13626 9881 13628
rect 9905 13626 9961 13628
rect 9665 13574 9691 13626
rect 9691 13574 9721 13626
rect 9745 13574 9755 13626
rect 9755 13574 9801 13626
rect 9825 13574 9871 13626
rect 9871 13574 9881 13626
rect 9905 13574 9935 13626
rect 9935 13574 9961 13626
rect 9665 13572 9721 13574
rect 9745 13572 9801 13574
rect 9825 13572 9881 13574
rect 9905 13572 9961 13574
rect 7488 13082 7544 13084
rect 7568 13082 7624 13084
rect 7648 13082 7704 13084
rect 7728 13082 7784 13084
rect 7488 13030 7514 13082
rect 7514 13030 7544 13082
rect 7568 13030 7578 13082
rect 7578 13030 7624 13082
rect 7648 13030 7694 13082
rect 7694 13030 7704 13082
rect 7728 13030 7758 13082
rect 7758 13030 7784 13082
rect 7488 13028 7544 13030
rect 7568 13028 7624 13030
rect 7648 13028 7704 13030
rect 7728 13028 7784 13030
rect 5310 12538 5366 12540
rect 5390 12538 5446 12540
rect 5470 12538 5526 12540
rect 5550 12538 5606 12540
rect 5310 12486 5336 12538
rect 5336 12486 5366 12538
rect 5390 12486 5400 12538
rect 5400 12486 5446 12538
rect 5470 12486 5516 12538
rect 5516 12486 5526 12538
rect 5550 12486 5580 12538
rect 5580 12486 5606 12538
rect 5310 12484 5366 12486
rect 5390 12484 5446 12486
rect 5470 12484 5526 12486
rect 5550 12484 5606 12486
rect 9665 12538 9721 12540
rect 9745 12538 9801 12540
rect 9825 12538 9881 12540
rect 9905 12538 9961 12540
rect 9665 12486 9691 12538
rect 9691 12486 9721 12538
rect 9745 12486 9755 12538
rect 9755 12486 9801 12538
rect 9825 12486 9871 12538
rect 9871 12486 9881 12538
rect 9905 12486 9935 12538
rect 9935 12486 9961 12538
rect 9665 12484 9721 12486
rect 9745 12484 9801 12486
rect 9825 12484 9881 12486
rect 9905 12484 9961 12486
rect 7488 11994 7544 11996
rect 7568 11994 7624 11996
rect 7648 11994 7704 11996
rect 7728 11994 7784 11996
rect 7488 11942 7514 11994
rect 7514 11942 7544 11994
rect 7568 11942 7578 11994
rect 7578 11942 7624 11994
rect 7648 11942 7694 11994
rect 7694 11942 7704 11994
rect 7728 11942 7758 11994
rect 7758 11942 7784 11994
rect 7488 11940 7544 11942
rect 7568 11940 7624 11942
rect 7648 11940 7704 11942
rect 7728 11940 7784 11942
rect 5310 11450 5366 11452
rect 5390 11450 5446 11452
rect 5470 11450 5526 11452
rect 5550 11450 5606 11452
rect 5310 11398 5336 11450
rect 5336 11398 5366 11450
rect 5390 11398 5400 11450
rect 5400 11398 5446 11450
rect 5470 11398 5516 11450
rect 5516 11398 5526 11450
rect 5550 11398 5580 11450
rect 5580 11398 5606 11450
rect 5310 11396 5366 11398
rect 5390 11396 5446 11398
rect 5470 11396 5526 11398
rect 5550 11396 5606 11398
rect 9665 11450 9721 11452
rect 9745 11450 9801 11452
rect 9825 11450 9881 11452
rect 9905 11450 9961 11452
rect 9665 11398 9691 11450
rect 9691 11398 9721 11450
rect 9745 11398 9755 11450
rect 9755 11398 9801 11450
rect 9825 11398 9871 11450
rect 9871 11398 9881 11450
rect 9905 11398 9935 11450
rect 9935 11398 9961 11450
rect 9665 11396 9721 11398
rect 9745 11396 9801 11398
rect 9825 11396 9881 11398
rect 9905 11396 9961 11398
rect 7488 10906 7544 10908
rect 7568 10906 7624 10908
rect 7648 10906 7704 10908
rect 7728 10906 7784 10908
rect 7488 10854 7514 10906
rect 7514 10854 7544 10906
rect 7568 10854 7578 10906
rect 7578 10854 7624 10906
rect 7648 10854 7694 10906
rect 7694 10854 7704 10906
rect 7728 10854 7758 10906
rect 7758 10854 7784 10906
rect 7488 10852 7544 10854
rect 7568 10852 7624 10854
rect 7648 10852 7704 10854
rect 7728 10852 7784 10854
rect 5310 10362 5366 10364
rect 5390 10362 5446 10364
rect 5470 10362 5526 10364
rect 5550 10362 5606 10364
rect 5310 10310 5336 10362
rect 5336 10310 5366 10362
rect 5390 10310 5400 10362
rect 5400 10310 5446 10362
rect 5470 10310 5516 10362
rect 5516 10310 5526 10362
rect 5550 10310 5580 10362
rect 5580 10310 5606 10362
rect 5310 10308 5366 10310
rect 5390 10308 5446 10310
rect 5470 10308 5526 10310
rect 5550 10308 5606 10310
rect 3133 9818 3189 9820
rect 3213 9818 3269 9820
rect 3293 9818 3349 9820
rect 3373 9818 3429 9820
rect 3133 9766 3159 9818
rect 3159 9766 3189 9818
rect 3213 9766 3223 9818
rect 3223 9766 3269 9818
rect 3293 9766 3339 9818
rect 3339 9766 3349 9818
rect 3373 9766 3403 9818
rect 3403 9766 3429 9818
rect 3133 9764 3189 9766
rect 3213 9764 3269 9766
rect 3293 9764 3349 9766
rect 3373 9764 3429 9766
rect 5310 9274 5366 9276
rect 5390 9274 5446 9276
rect 5470 9274 5526 9276
rect 5550 9274 5606 9276
rect 5310 9222 5336 9274
rect 5336 9222 5366 9274
rect 5390 9222 5400 9274
rect 5400 9222 5446 9274
rect 5470 9222 5516 9274
rect 5516 9222 5526 9274
rect 5550 9222 5580 9274
rect 5580 9222 5606 9274
rect 5310 9220 5366 9222
rect 5390 9220 5446 9222
rect 5470 9220 5526 9222
rect 5550 9220 5606 9222
rect 7488 9818 7544 9820
rect 7568 9818 7624 9820
rect 7648 9818 7704 9820
rect 7728 9818 7784 9820
rect 7488 9766 7514 9818
rect 7514 9766 7544 9818
rect 7568 9766 7578 9818
rect 7578 9766 7624 9818
rect 7648 9766 7694 9818
rect 7694 9766 7704 9818
rect 7728 9766 7758 9818
rect 7758 9766 7784 9818
rect 7488 9764 7544 9766
rect 7568 9764 7624 9766
rect 7648 9764 7704 9766
rect 7728 9764 7784 9766
rect 3133 8730 3189 8732
rect 3213 8730 3269 8732
rect 3293 8730 3349 8732
rect 3373 8730 3429 8732
rect 3133 8678 3159 8730
rect 3159 8678 3189 8730
rect 3213 8678 3223 8730
rect 3223 8678 3269 8730
rect 3293 8678 3339 8730
rect 3339 8678 3349 8730
rect 3373 8678 3403 8730
rect 3403 8678 3429 8730
rect 3133 8676 3189 8678
rect 3213 8676 3269 8678
rect 3293 8676 3349 8678
rect 3373 8676 3429 8678
rect 7488 8730 7544 8732
rect 7568 8730 7624 8732
rect 7648 8730 7704 8732
rect 7728 8730 7784 8732
rect 7488 8678 7514 8730
rect 7514 8678 7544 8730
rect 7568 8678 7578 8730
rect 7578 8678 7624 8730
rect 7648 8678 7694 8730
rect 7694 8678 7704 8730
rect 7728 8678 7758 8730
rect 7758 8678 7784 8730
rect 7488 8676 7544 8678
rect 7568 8676 7624 8678
rect 7648 8676 7704 8678
rect 7728 8676 7784 8678
rect 5310 8186 5366 8188
rect 5390 8186 5446 8188
rect 5470 8186 5526 8188
rect 5550 8186 5606 8188
rect 5310 8134 5336 8186
rect 5336 8134 5366 8186
rect 5390 8134 5400 8186
rect 5400 8134 5446 8186
rect 5470 8134 5516 8186
rect 5516 8134 5526 8186
rect 5550 8134 5580 8186
rect 5580 8134 5606 8186
rect 5310 8132 5366 8134
rect 5390 8132 5446 8134
rect 5470 8132 5526 8134
rect 5550 8132 5606 8134
rect 3133 7642 3189 7644
rect 3213 7642 3269 7644
rect 3293 7642 3349 7644
rect 3373 7642 3429 7644
rect 3133 7590 3159 7642
rect 3159 7590 3189 7642
rect 3213 7590 3223 7642
rect 3223 7590 3269 7642
rect 3293 7590 3339 7642
rect 3339 7590 3349 7642
rect 3373 7590 3403 7642
rect 3403 7590 3429 7642
rect 3133 7588 3189 7590
rect 3213 7588 3269 7590
rect 3293 7588 3349 7590
rect 3373 7588 3429 7590
rect 7488 7642 7544 7644
rect 7568 7642 7624 7644
rect 7648 7642 7704 7644
rect 7728 7642 7784 7644
rect 7488 7590 7514 7642
rect 7514 7590 7544 7642
rect 7568 7590 7578 7642
rect 7578 7590 7624 7642
rect 7648 7590 7694 7642
rect 7694 7590 7704 7642
rect 7728 7590 7758 7642
rect 7758 7590 7784 7642
rect 7488 7588 7544 7590
rect 7568 7588 7624 7590
rect 7648 7588 7704 7590
rect 7728 7588 7784 7590
rect 5310 7098 5366 7100
rect 5390 7098 5446 7100
rect 5470 7098 5526 7100
rect 5550 7098 5606 7100
rect 5310 7046 5336 7098
rect 5336 7046 5366 7098
rect 5390 7046 5400 7098
rect 5400 7046 5446 7098
rect 5470 7046 5516 7098
rect 5516 7046 5526 7098
rect 5550 7046 5580 7098
rect 5580 7046 5606 7098
rect 5310 7044 5366 7046
rect 5390 7044 5446 7046
rect 5470 7044 5526 7046
rect 5550 7044 5606 7046
rect 3133 6554 3189 6556
rect 3213 6554 3269 6556
rect 3293 6554 3349 6556
rect 3373 6554 3429 6556
rect 3133 6502 3159 6554
rect 3159 6502 3189 6554
rect 3213 6502 3223 6554
rect 3223 6502 3269 6554
rect 3293 6502 3339 6554
rect 3339 6502 3349 6554
rect 3373 6502 3403 6554
rect 3403 6502 3429 6554
rect 3133 6500 3189 6502
rect 3213 6500 3269 6502
rect 3293 6500 3349 6502
rect 3373 6500 3429 6502
rect 7488 6554 7544 6556
rect 7568 6554 7624 6556
rect 7648 6554 7704 6556
rect 7728 6554 7784 6556
rect 7488 6502 7514 6554
rect 7514 6502 7544 6554
rect 7568 6502 7578 6554
rect 7578 6502 7624 6554
rect 7648 6502 7694 6554
rect 7694 6502 7704 6554
rect 7728 6502 7758 6554
rect 7758 6502 7784 6554
rect 7488 6500 7544 6502
rect 7568 6500 7624 6502
rect 7648 6500 7704 6502
rect 7728 6500 7784 6502
rect 5310 6010 5366 6012
rect 5390 6010 5446 6012
rect 5470 6010 5526 6012
rect 5550 6010 5606 6012
rect 5310 5958 5336 6010
rect 5336 5958 5366 6010
rect 5390 5958 5400 6010
rect 5400 5958 5446 6010
rect 5470 5958 5516 6010
rect 5516 5958 5526 6010
rect 5550 5958 5580 6010
rect 5580 5958 5606 6010
rect 5310 5956 5366 5958
rect 5390 5956 5446 5958
rect 5470 5956 5526 5958
rect 5550 5956 5606 5958
rect 3133 5466 3189 5468
rect 3213 5466 3269 5468
rect 3293 5466 3349 5468
rect 3373 5466 3429 5468
rect 3133 5414 3159 5466
rect 3159 5414 3189 5466
rect 3213 5414 3223 5466
rect 3223 5414 3269 5466
rect 3293 5414 3339 5466
rect 3339 5414 3349 5466
rect 3373 5414 3403 5466
rect 3403 5414 3429 5466
rect 3133 5412 3189 5414
rect 3213 5412 3269 5414
rect 3293 5412 3349 5414
rect 3373 5412 3429 5414
rect 7488 5466 7544 5468
rect 7568 5466 7624 5468
rect 7648 5466 7704 5468
rect 7728 5466 7784 5468
rect 7488 5414 7514 5466
rect 7514 5414 7544 5466
rect 7568 5414 7578 5466
rect 7578 5414 7624 5466
rect 7648 5414 7694 5466
rect 7694 5414 7704 5466
rect 7728 5414 7758 5466
rect 7758 5414 7784 5466
rect 7488 5412 7544 5414
rect 7568 5412 7624 5414
rect 7648 5412 7704 5414
rect 7728 5412 7784 5414
rect 5310 4922 5366 4924
rect 5390 4922 5446 4924
rect 5470 4922 5526 4924
rect 5550 4922 5606 4924
rect 5310 4870 5336 4922
rect 5336 4870 5366 4922
rect 5390 4870 5400 4922
rect 5400 4870 5446 4922
rect 5470 4870 5516 4922
rect 5516 4870 5526 4922
rect 5550 4870 5580 4922
rect 5580 4870 5606 4922
rect 5310 4868 5366 4870
rect 5390 4868 5446 4870
rect 5470 4868 5526 4870
rect 5550 4868 5606 4870
rect 3133 4378 3189 4380
rect 3213 4378 3269 4380
rect 3293 4378 3349 4380
rect 3373 4378 3429 4380
rect 3133 4326 3159 4378
rect 3159 4326 3189 4378
rect 3213 4326 3223 4378
rect 3223 4326 3269 4378
rect 3293 4326 3339 4378
rect 3339 4326 3349 4378
rect 3373 4326 3403 4378
rect 3403 4326 3429 4378
rect 3133 4324 3189 4326
rect 3213 4324 3269 4326
rect 3293 4324 3349 4326
rect 3373 4324 3429 4326
rect 7488 4378 7544 4380
rect 7568 4378 7624 4380
rect 7648 4378 7704 4380
rect 7728 4378 7784 4380
rect 7488 4326 7514 4378
rect 7514 4326 7544 4378
rect 7568 4326 7578 4378
rect 7578 4326 7624 4378
rect 7648 4326 7694 4378
rect 7694 4326 7704 4378
rect 7728 4326 7758 4378
rect 7758 4326 7784 4378
rect 7488 4324 7544 4326
rect 7568 4324 7624 4326
rect 7648 4324 7704 4326
rect 7728 4324 7784 4326
rect 5310 3834 5366 3836
rect 5390 3834 5446 3836
rect 5470 3834 5526 3836
rect 5550 3834 5606 3836
rect 5310 3782 5336 3834
rect 5336 3782 5366 3834
rect 5390 3782 5400 3834
rect 5400 3782 5446 3834
rect 5470 3782 5516 3834
rect 5516 3782 5526 3834
rect 5550 3782 5580 3834
rect 5580 3782 5606 3834
rect 5310 3780 5366 3782
rect 5390 3780 5446 3782
rect 5470 3780 5526 3782
rect 5550 3780 5606 3782
rect 3133 3290 3189 3292
rect 3213 3290 3269 3292
rect 3293 3290 3349 3292
rect 3373 3290 3429 3292
rect 3133 3238 3159 3290
rect 3159 3238 3189 3290
rect 3213 3238 3223 3290
rect 3223 3238 3269 3290
rect 3293 3238 3339 3290
rect 3339 3238 3349 3290
rect 3373 3238 3403 3290
rect 3403 3238 3429 3290
rect 3133 3236 3189 3238
rect 3213 3236 3269 3238
rect 3293 3236 3349 3238
rect 3373 3236 3429 3238
rect 7488 3290 7544 3292
rect 7568 3290 7624 3292
rect 7648 3290 7704 3292
rect 7728 3290 7784 3292
rect 7488 3238 7514 3290
rect 7514 3238 7544 3290
rect 7568 3238 7578 3290
rect 7578 3238 7624 3290
rect 7648 3238 7694 3290
rect 7694 3238 7704 3290
rect 7728 3238 7758 3290
rect 7758 3238 7784 3290
rect 7488 3236 7544 3238
rect 7568 3236 7624 3238
rect 7648 3236 7704 3238
rect 7728 3236 7784 3238
rect 5310 2746 5366 2748
rect 5390 2746 5446 2748
rect 5470 2746 5526 2748
rect 5550 2746 5606 2748
rect 5310 2694 5336 2746
rect 5336 2694 5366 2746
rect 5390 2694 5400 2746
rect 5400 2694 5446 2746
rect 5470 2694 5516 2746
rect 5516 2694 5526 2746
rect 5550 2694 5580 2746
rect 5580 2694 5606 2746
rect 5310 2692 5366 2694
rect 5390 2692 5446 2694
rect 5470 2692 5526 2694
rect 5550 2692 5606 2694
rect 9665 10362 9721 10364
rect 9745 10362 9801 10364
rect 9825 10362 9881 10364
rect 9905 10362 9961 10364
rect 9665 10310 9691 10362
rect 9691 10310 9721 10362
rect 9745 10310 9755 10362
rect 9755 10310 9801 10362
rect 9825 10310 9871 10362
rect 9871 10310 9881 10362
rect 9905 10310 9935 10362
rect 9935 10310 9961 10362
rect 9665 10308 9721 10310
rect 9745 10308 9801 10310
rect 9825 10308 9881 10310
rect 9905 10308 9961 10310
rect 9665 9274 9721 9276
rect 9745 9274 9801 9276
rect 9825 9274 9881 9276
rect 9905 9274 9961 9276
rect 9665 9222 9691 9274
rect 9691 9222 9721 9274
rect 9745 9222 9755 9274
rect 9755 9222 9801 9274
rect 9825 9222 9871 9274
rect 9871 9222 9881 9274
rect 9905 9222 9935 9274
rect 9935 9222 9961 9274
rect 9665 9220 9721 9222
rect 9745 9220 9801 9222
rect 9825 9220 9881 9222
rect 9905 9220 9961 9222
rect 9665 8186 9721 8188
rect 9745 8186 9801 8188
rect 9825 8186 9881 8188
rect 9905 8186 9961 8188
rect 9665 8134 9691 8186
rect 9691 8134 9721 8186
rect 9745 8134 9755 8186
rect 9755 8134 9801 8186
rect 9825 8134 9871 8186
rect 9871 8134 9881 8186
rect 9905 8134 9935 8186
rect 9935 8134 9961 8186
rect 9665 8132 9721 8134
rect 9745 8132 9801 8134
rect 9825 8132 9881 8134
rect 9905 8132 9961 8134
rect 9665 7098 9721 7100
rect 9745 7098 9801 7100
rect 9825 7098 9881 7100
rect 9905 7098 9961 7100
rect 9665 7046 9691 7098
rect 9691 7046 9721 7098
rect 9745 7046 9755 7098
rect 9755 7046 9801 7098
rect 9825 7046 9871 7098
rect 9871 7046 9881 7098
rect 9905 7046 9935 7098
rect 9935 7046 9961 7098
rect 9665 7044 9721 7046
rect 9745 7044 9801 7046
rect 9825 7044 9881 7046
rect 9905 7044 9961 7046
rect 9665 6010 9721 6012
rect 9745 6010 9801 6012
rect 9825 6010 9881 6012
rect 9905 6010 9961 6012
rect 9665 5958 9691 6010
rect 9691 5958 9721 6010
rect 9745 5958 9755 6010
rect 9755 5958 9801 6010
rect 9825 5958 9871 6010
rect 9871 5958 9881 6010
rect 9905 5958 9935 6010
rect 9935 5958 9961 6010
rect 9665 5956 9721 5958
rect 9745 5956 9801 5958
rect 9825 5956 9881 5958
rect 9905 5956 9961 5958
rect 9665 4922 9721 4924
rect 9745 4922 9801 4924
rect 9825 4922 9881 4924
rect 9905 4922 9961 4924
rect 9665 4870 9691 4922
rect 9691 4870 9721 4922
rect 9745 4870 9755 4922
rect 9755 4870 9801 4922
rect 9825 4870 9871 4922
rect 9871 4870 9881 4922
rect 9905 4870 9935 4922
rect 9935 4870 9961 4922
rect 9665 4868 9721 4870
rect 9745 4868 9801 4870
rect 9825 4868 9881 4870
rect 9905 4868 9961 4870
rect 9665 3834 9721 3836
rect 9745 3834 9801 3836
rect 9825 3834 9881 3836
rect 9905 3834 9961 3836
rect 9665 3782 9691 3834
rect 9691 3782 9721 3834
rect 9745 3782 9755 3834
rect 9755 3782 9801 3834
rect 9825 3782 9871 3834
rect 9871 3782 9881 3834
rect 9905 3782 9935 3834
rect 9935 3782 9961 3834
rect 9665 3780 9721 3782
rect 9745 3780 9801 3782
rect 9825 3780 9881 3782
rect 9905 3780 9961 3782
rect 11842 15258 11898 15260
rect 11922 15258 11978 15260
rect 12002 15258 12058 15260
rect 12082 15258 12138 15260
rect 11842 15206 11868 15258
rect 11868 15206 11898 15258
rect 11922 15206 11932 15258
rect 11932 15206 11978 15258
rect 12002 15206 12048 15258
rect 12048 15206 12058 15258
rect 12082 15206 12112 15258
rect 12112 15206 12138 15258
rect 11842 15204 11898 15206
rect 11922 15204 11978 15206
rect 12002 15204 12058 15206
rect 12082 15204 12138 15206
rect 11842 14170 11898 14172
rect 11922 14170 11978 14172
rect 12002 14170 12058 14172
rect 12082 14170 12138 14172
rect 11842 14118 11868 14170
rect 11868 14118 11898 14170
rect 11922 14118 11932 14170
rect 11932 14118 11978 14170
rect 12002 14118 12048 14170
rect 12048 14118 12058 14170
rect 12082 14118 12112 14170
rect 12112 14118 12138 14170
rect 11842 14116 11898 14118
rect 11922 14116 11978 14118
rect 12002 14116 12058 14118
rect 12082 14116 12138 14118
rect 11842 13082 11898 13084
rect 11922 13082 11978 13084
rect 12002 13082 12058 13084
rect 12082 13082 12138 13084
rect 11842 13030 11868 13082
rect 11868 13030 11898 13082
rect 11922 13030 11932 13082
rect 11932 13030 11978 13082
rect 12002 13030 12048 13082
rect 12048 13030 12058 13082
rect 12082 13030 12112 13082
rect 12112 13030 12138 13082
rect 11842 13028 11898 13030
rect 11922 13028 11978 13030
rect 12002 13028 12058 13030
rect 12082 13028 12138 13030
rect 11842 11994 11898 11996
rect 11922 11994 11978 11996
rect 12002 11994 12058 11996
rect 12082 11994 12138 11996
rect 11842 11942 11868 11994
rect 11868 11942 11898 11994
rect 11922 11942 11932 11994
rect 11932 11942 11978 11994
rect 12002 11942 12048 11994
rect 12048 11942 12058 11994
rect 12082 11942 12112 11994
rect 12112 11942 12138 11994
rect 11842 11940 11898 11942
rect 11922 11940 11978 11942
rect 12002 11940 12058 11942
rect 12082 11940 12138 11942
rect 13450 11620 13506 11656
rect 13450 11600 13452 11620
rect 13452 11600 13504 11620
rect 13504 11600 13506 11620
rect 11842 10906 11898 10908
rect 11922 10906 11978 10908
rect 12002 10906 12058 10908
rect 12082 10906 12138 10908
rect 11842 10854 11868 10906
rect 11868 10854 11898 10906
rect 11922 10854 11932 10906
rect 11932 10854 11978 10906
rect 12002 10854 12048 10906
rect 12048 10854 12058 10906
rect 12082 10854 12112 10906
rect 12112 10854 12138 10906
rect 11842 10852 11898 10854
rect 11922 10852 11978 10854
rect 12002 10852 12058 10854
rect 12082 10852 12138 10854
rect 11842 9818 11898 9820
rect 11922 9818 11978 9820
rect 12002 9818 12058 9820
rect 12082 9818 12138 9820
rect 11842 9766 11868 9818
rect 11868 9766 11898 9818
rect 11922 9766 11932 9818
rect 11932 9766 11978 9818
rect 12002 9766 12048 9818
rect 12048 9766 12058 9818
rect 12082 9766 12112 9818
rect 12112 9766 12138 9818
rect 11842 9764 11898 9766
rect 11922 9764 11978 9766
rect 12002 9764 12058 9766
rect 12082 9764 12138 9766
rect 11842 8730 11898 8732
rect 11922 8730 11978 8732
rect 12002 8730 12058 8732
rect 12082 8730 12138 8732
rect 11842 8678 11868 8730
rect 11868 8678 11898 8730
rect 11922 8678 11932 8730
rect 11932 8678 11978 8730
rect 12002 8678 12048 8730
rect 12048 8678 12058 8730
rect 12082 8678 12112 8730
rect 12112 8678 12138 8730
rect 11842 8676 11898 8678
rect 11922 8676 11978 8678
rect 12002 8676 12058 8678
rect 12082 8676 12138 8678
rect 11842 7642 11898 7644
rect 11922 7642 11978 7644
rect 12002 7642 12058 7644
rect 12082 7642 12138 7644
rect 11842 7590 11868 7642
rect 11868 7590 11898 7642
rect 11922 7590 11932 7642
rect 11932 7590 11978 7642
rect 12002 7590 12048 7642
rect 12048 7590 12058 7642
rect 12082 7590 12112 7642
rect 12112 7590 12138 7642
rect 11842 7588 11898 7590
rect 11922 7588 11978 7590
rect 12002 7588 12058 7590
rect 12082 7588 12138 7590
rect 11842 6554 11898 6556
rect 11922 6554 11978 6556
rect 12002 6554 12058 6556
rect 12082 6554 12138 6556
rect 11842 6502 11868 6554
rect 11868 6502 11898 6554
rect 11922 6502 11932 6554
rect 11932 6502 11978 6554
rect 12002 6502 12048 6554
rect 12048 6502 12058 6554
rect 12082 6502 12112 6554
rect 12112 6502 12138 6554
rect 11842 6500 11898 6502
rect 11922 6500 11978 6502
rect 12002 6500 12058 6502
rect 12082 6500 12138 6502
rect 11842 5466 11898 5468
rect 11922 5466 11978 5468
rect 12002 5466 12058 5468
rect 12082 5466 12138 5468
rect 11842 5414 11868 5466
rect 11868 5414 11898 5466
rect 11922 5414 11932 5466
rect 11932 5414 11978 5466
rect 12002 5414 12048 5466
rect 12048 5414 12058 5466
rect 12082 5414 12112 5466
rect 12112 5414 12138 5466
rect 11842 5412 11898 5414
rect 11922 5412 11978 5414
rect 12002 5412 12058 5414
rect 12082 5412 12138 5414
rect 11842 4378 11898 4380
rect 11922 4378 11978 4380
rect 12002 4378 12058 4380
rect 12082 4378 12138 4380
rect 11842 4326 11868 4378
rect 11868 4326 11898 4378
rect 11922 4326 11932 4378
rect 11932 4326 11978 4378
rect 12002 4326 12048 4378
rect 12048 4326 12058 4378
rect 12082 4326 12112 4378
rect 12112 4326 12138 4378
rect 11842 4324 11898 4326
rect 11922 4324 11978 4326
rect 12002 4324 12058 4326
rect 12082 4324 12138 4326
rect 11842 3290 11898 3292
rect 11922 3290 11978 3292
rect 12002 3290 12058 3292
rect 12082 3290 12138 3292
rect 11842 3238 11868 3290
rect 11868 3238 11898 3290
rect 11922 3238 11932 3290
rect 11932 3238 11978 3290
rect 12002 3238 12048 3290
rect 12048 3238 12058 3290
rect 12082 3238 12112 3290
rect 12112 3238 12138 3290
rect 11842 3236 11898 3238
rect 11922 3236 11978 3238
rect 12002 3236 12058 3238
rect 12082 3236 12138 3238
rect 9665 2746 9721 2748
rect 9745 2746 9801 2748
rect 9825 2746 9881 2748
rect 9905 2746 9961 2748
rect 9665 2694 9691 2746
rect 9691 2694 9721 2746
rect 9745 2694 9755 2746
rect 9755 2694 9801 2746
rect 9825 2694 9871 2746
rect 9871 2694 9881 2746
rect 9905 2694 9935 2746
rect 9935 2694 9961 2746
rect 9665 2692 9721 2694
rect 9745 2692 9801 2694
rect 9825 2692 9881 2694
rect 9905 2692 9961 2694
rect 3133 2202 3189 2204
rect 3213 2202 3269 2204
rect 3293 2202 3349 2204
rect 3373 2202 3429 2204
rect 3133 2150 3159 2202
rect 3159 2150 3189 2202
rect 3213 2150 3223 2202
rect 3223 2150 3269 2202
rect 3293 2150 3339 2202
rect 3339 2150 3349 2202
rect 3373 2150 3403 2202
rect 3403 2150 3429 2202
rect 3133 2148 3189 2150
rect 3213 2148 3269 2150
rect 3293 2148 3349 2150
rect 3373 2148 3429 2150
rect 7488 2202 7544 2204
rect 7568 2202 7624 2204
rect 7648 2202 7704 2204
rect 7728 2202 7784 2204
rect 7488 2150 7514 2202
rect 7514 2150 7544 2202
rect 7568 2150 7578 2202
rect 7578 2150 7624 2202
rect 7648 2150 7694 2202
rect 7694 2150 7704 2202
rect 7728 2150 7758 2202
rect 7758 2150 7784 2202
rect 7488 2148 7544 2150
rect 7568 2148 7624 2150
rect 7648 2148 7704 2150
rect 7728 2148 7784 2150
rect 11842 2202 11898 2204
rect 11922 2202 11978 2204
rect 12002 2202 12058 2204
rect 12082 2202 12138 2204
rect 11842 2150 11868 2202
rect 11868 2150 11898 2202
rect 11922 2150 11932 2202
rect 11932 2150 11978 2202
rect 12002 2150 12048 2202
rect 12048 2150 12058 2202
rect 12082 2150 12112 2202
rect 12112 2150 12138 2202
rect 11842 2148 11898 2150
rect 11922 2148 11978 2150
rect 12002 2148 12058 2150
rect 12082 2148 12138 2150
rect 13450 720 13506 776
<< metal3 >>
rect 3121 15264 3441 15265
rect 3121 15200 3129 15264
rect 3193 15200 3209 15264
rect 3273 15200 3289 15264
rect 3353 15200 3369 15264
rect 3433 15200 3441 15264
rect 3121 15199 3441 15200
rect 7476 15264 7796 15265
rect 7476 15200 7484 15264
rect 7548 15200 7564 15264
rect 7628 15200 7644 15264
rect 7708 15200 7724 15264
rect 7788 15200 7796 15264
rect 7476 15199 7796 15200
rect 11830 15264 12150 15265
rect 11830 15200 11838 15264
rect 11902 15200 11918 15264
rect 11982 15200 11998 15264
rect 12062 15200 12078 15264
rect 12142 15200 12150 15264
rect 11830 15199 12150 15200
rect 5298 14720 5618 14721
rect 5298 14656 5306 14720
rect 5370 14656 5386 14720
rect 5450 14656 5466 14720
rect 5530 14656 5546 14720
rect 5610 14656 5618 14720
rect 5298 14655 5618 14656
rect 9653 14720 9973 14721
rect 9653 14656 9661 14720
rect 9725 14656 9741 14720
rect 9805 14656 9821 14720
rect 9885 14656 9901 14720
rect 9965 14656 9973 14720
rect 9653 14655 9973 14656
rect 3121 14176 3441 14177
rect 3121 14112 3129 14176
rect 3193 14112 3209 14176
rect 3273 14112 3289 14176
rect 3353 14112 3369 14176
rect 3433 14112 3441 14176
rect 3121 14111 3441 14112
rect 7476 14176 7796 14177
rect 7476 14112 7484 14176
rect 7548 14112 7564 14176
rect 7628 14112 7644 14176
rect 7708 14112 7724 14176
rect 7788 14112 7796 14176
rect 7476 14111 7796 14112
rect 11830 14176 12150 14177
rect 11830 14112 11838 14176
rect 11902 14112 11918 14176
rect 11982 14112 11998 14176
rect 12062 14112 12078 14176
rect 12142 14112 12150 14176
rect 11830 14111 12150 14112
rect 5298 13632 5618 13633
rect 5298 13568 5306 13632
rect 5370 13568 5386 13632
rect 5450 13568 5466 13632
rect 5530 13568 5546 13632
rect 5610 13568 5618 13632
rect 5298 13567 5618 13568
rect 9653 13632 9973 13633
rect 9653 13568 9661 13632
rect 9725 13568 9741 13632
rect 9805 13568 9821 13632
rect 9885 13568 9901 13632
rect 9965 13568 9973 13632
rect 9653 13567 9973 13568
rect 3121 13088 3441 13089
rect 3121 13024 3129 13088
rect 3193 13024 3209 13088
rect 3273 13024 3289 13088
rect 3353 13024 3369 13088
rect 3433 13024 3441 13088
rect 3121 13023 3441 13024
rect 7476 13088 7796 13089
rect 7476 13024 7484 13088
rect 7548 13024 7564 13088
rect 7628 13024 7644 13088
rect 7708 13024 7724 13088
rect 7788 13024 7796 13088
rect 7476 13023 7796 13024
rect 11830 13088 12150 13089
rect 11830 13024 11838 13088
rect 11902 13024 11918 13088
rect 11982 13024 11998 13088
rect 12062 13024 12078 13088
rect 12142 13024 12150 13088
rect 11830 13023 12150 13024
rect 5298 12544 5618 12545
rect 5298 12480 5306 12544
rect 5370 12480 5386 12544
rect 5450 12480 5466 12544
rect 5530 12480 5546 12544
rect 5610 12480 5618 12544
rect 5298 12479 5618 12480
rect 9653 12544 9973 12545
rect 9653 12480 9661 12544
rect 9725 12480 9741 12544
rect 9805 12480 9821 12544
rect 9885 12480 9901 12544
rect 9965 12480 9973 12544
rect 9653 12479 9973 12480
rect 3121 12000 3441 12001
rect 3121 11936 3129 12000
rect 3193 11936 3209 12000
rect 3273 11936 3289 12000
rect 3353 11936 3369 12000
rect 3433 11936 3441 12000
rect 3121 11935 3441 11936
rect 7476 12000 7796 12001
rect 7476 11936 7484 12000
rect 7548 11936 7564 12000
rect 7628 11936 7644 12000
rect 7708 11936 7724 12000
rect 7788 11936 7796 12000
rect 7476 11935 7796 11936
rect 11830 12000 12150 12001
rect 11830 11936 11838 12000
rect 11902 11936 11918 12000
rect 11982 11936 11998 12000
rect 12062 11936 12078 12000
rect 12142 11936 12150 12000
rect 11830 11935 12150 11936
rect 13445 11658 13511 11661
rect 14491 11658 15291 11688
rect 13445 11656 15291 11658
rect 13445 11600 13450 11656
rect 13506 11600 15291 11656
rect 13445 11598 15291 11600
rect 13445 11595 13511 11598
rect 14491 11568 15291 11598
rect 5298 11456 5618 11457
rect 5298 11392 5306 11456
rect 5370 11392 5386 11456
rect 5450 11392 5466 11456
rect 5530 11392 5546 11456
rect 5610 11392 5618 11456
rect 5298 11391 5618 11392
rect 9653 11456 9973 11457
rect 9653 11392 9661 11456
rect 9725 11392 9741 11456
rect 9805 11392 9821 11456
rect 9885 11392 9901 11456
rect 9965 11392 9973 11456
rect 9653 11391 9973 11392
rect 0 10978 800 11008
rect 1761 10978 1827 10981
rect 0 10976 1827 10978
rect 0 10920 1766 10976
rect 1822 10920 1827 10976
rect 0 10918 1827 10920
rect 0 10888 800 10918
rect 1761 10915 1827 10918
rect 3121 10912 3441 10913
rect 3121 10848 3129 10912
rect 3193 10848 3209 10912
rect 3273 10848 3289 10912
rect 3353 10848 3369 10912
rect 3433 10848 3441 10912
rect 3121 10847 3441 10848
rect 7476 10912 7796 10913
rect 7476 10848 7484 10912
rect 7548 10848 7564 10912
rect 7628 10848 7644 10912
rect 7708 10848 7724 10912
rect 7788 10848 7796 10912
rect 7476 10847 7796 10848
rect 11830 10912 12150 10913
rect 11830 10848 11838 10912
rect 11902 10848 11918 10912
rect 11982 10848 11998 10912
rect 12062 10848 12078 10912
rect 12142 10848 12150 10912
rect 11830 10847 12150 10848
rect 5298 10368 5618 10369
rect 5298 10304 5306 10368
rect 5370 10304 5386 10368
rect 5450 10304 5466 10368
rect 5530 10304 5546 10368
rect 5610 10304 5618 10368
rect 5298 10303 5618 10304
rect 9653 10368 9973 10369
rect 9653 10304 9661 10368
rect 9725 10304 9741 10368
rect 9805 10304 9821 10368
rect 9885 10304 9901 10368
rect 9965 10304 9973 10368
rect 9653 10303 9973 10304
rect 3121 9824 3441 9825
rect 3121 9760 3129 9824
rect 3193 9760 3209 9824
rect 3273 9760 3289 9824
rect 3353 9760 3369 9824
rect 3433 9760 3441 9824
rect 3121 9759 3441 9760
rect 7476 9824 7796 9825
rect 7476 9760 7484 9824
rect 7548 9760 7564 9824
rect 7628 9760 7644 9824
rect 7708 9760 7724 9824
rect 7788 9760 7796 9824
rect 7476 9759 7796 9760
rect 11830 9824 12150 9825
rect 11830 9760 11838 9824
rect 11902 9760 11918 9824
rect 11982 9760 11998 9824
rect 12062 9760 12078 9824
rect 12142 9760 12150 9824
rect 11830 9759 12150 9760
rect 5298 9280 5618 9281
rect 5298 9216 5306 9280
rect 5370 9216 5386 9280
rect 5450 9216 5466 9280
rect 5530 9216 5546 9280
rect 5610 9216 5618 9280
rect 5298 9215 5618 9216
rect 9653 9280 9973 9281
rect 9653 9216 9661 9280
rect 9725 9216 9741 9280
rect 9805 9216 9821 9280
rect 9885 9216 9901 9280
rect 9965 9216 9973 9280
rect 9653 9215 9973 9216
rect 3121 8736 3441 8737
rect 3121 8672 3129 8736
rect 3193 8672 3209 8736
rect 3273 8672 3289 8736
rect 3353 8672 3369 8736
rect 3433 8672 3441 8736
rect 3121 8671 3441 8672
rect 7476 8736 7796 8737
rect 7476 8672 7484 8736
rect 7548 8672 7564 8736
rect 7628 8672 7644 8736
rect 7708 8672 7724 8736
rect 7788 8672 7796 8736
rect 7476 8671 7796 8672
rect 11830 8736 12150 8737
rect 11830 8672 11838 8736
rect 11902 8672 11918 8736
rect 11982 8672 11998 8736
rect 12062 8672 12078 8736
rect 12142 8672 12150 8736
rect 11830 8671 12150 8672
rect 5298 8192 5618 8193
rect 5298 8128 5306 8192
rect 5370 8128 5386 8192
rect 5450 8128 5466 8192
rect 5530 8128 5546 8192
rect 5610 8128 5618 8192
rect 5298 8127 5618 8128
rect 9653 8192 9973 8193
rect 9653 8128 9661 8192
rect 9725 8128 9741 8192
rect 9805 8128 9821 8192
rect 9885 8128 9901 8192
rect 9965 8128 9973 8192
rect 9653 8127 9973 8128
rect 3121 7648 3441 7649
rect 3121 7584 3129 7648
rect 3193 7584 3209 7648
rect 3273 7584 3289 7648
rect 3353 7584 3369 7648
rect 3433 7584 3441 7648
rect 3121 7583 3441 7584
rect 7476 7648 7796 7649
rect 7476 7584 7484 7648
rect 7548 7584 7564 7648
rect 7628 7584 7644 7648
rect 7708 7584 7724 7648
rect 7788 7584 7796 7648
rect 7476 7583 7796 7584
rect 11830 7648 12150 7649
rect 11830 7584 11838 7648
rect 11902 7584 11918 7648
rect 11982 7584 11998 7648
rect 12062 7584 12078 7648
rect 12142 7584 12150 7648
rect 11830 7583 12150 7584
rect 5298 7104 5618 7105
rect 5298 7040 5306 7104
rect 5370 7040 5386 7104
rect 5450 7040 5466 7104
rect 5530 7040 5546 7104
rect 5610 7040 5618 7104
rect 5298 7039 5618 7040
rect 9653 7104 9973 7105
rect 9653 7040 9661 7104
rect 9725 7040 9741 7104
rect 9805 7040 9821 7104
rect 9885 7040 9901 7104
rect 9965 7040 9973 7104
rect 9653 7039 9973 7040
rect 3121 6560 3441 6561
rect 3121 6496 3129 6560
rect 3193 6496 3209 6560
rect 3273 6496 3289 6560
rect 3353 6496 3369 6560
rect 3433 6496 3441 6560
rect 3121 6495 3441 6496
rect 7476 6560 7796 6561
rect 7476 6496 7484 6560
rect 7548 6496 7564 6560
rect 7628 6496 7644 6560
rect 7708 6496 7724 6560
rect 7788 6496 7796 6560
rect 7476 6495 7796 6496
rect 11830 6560 12150 6561
rect 11830 6496 11838 6560
rect 11902 6496 11918 6560
rect 11982 6496 11998 6560
rect 12062 6496 12078 6560
rect 12142 6496 12150 6560
rect 11830 6495 12150 6496
rect 5298 6016 5618 6017
rect 5298 5952 5306 6016
rect 5370 5952 5386 6016
rect 5450 5952 5466 6016
rect 5530 5952 5546 6016
rect 5610 5952 5618 6016
rect 5298 5951 5618 5952
rect 9653 6016 9973 6017
rect 9653 5952 9661 6016
rect 9725 5952 9741 6016
rect 9805 5952 9821 6016
rect 9885 5952 9901 6016
rect 9965 5952 9973 6016
rect 9653 5951 9973 5952
rect 3121 5472 3441 5473
rect 3121 5408 3129 5472
rect 3193 5408 3209 5472
rect 3273 5408 3289 5472
rect 3353 5408 3369 5472
rect 3433 5408 3441 5472
rect 3121 5407 3441 5408
rect 7476 5472 7796 5473
rect 7476 5408 7484 5472
rect 7548 5408 7564 5472
rect 7628 5408 7644 5472
rect 7708 5408 7724 5472
rect 7788 5408 7796 5472
rect 7476 5407 7796 5408
rect 11830 5472 12150 5473
rect 11830 5408 11838 5472
rect 11902 5408 11918 5472
rect 11982 5408 11998 5472
rect 12062 5408 12078 5472
rect 12142 5408 12150 5472
rect 11830 5407 12150 5408
rect 5298 4928 5618 4929
rect 5298 4864 5306 4928
rect 5370 4864 5386 4928
rect 5450 4864 5466 4928
rect 5530 4864 5546 4928
rect 5610 4864 5618 4928
rect 5298 4863 5618 4864
rect 9653 4928 9973 4929
rect 9653 4864 9661 4928
rect 9725 4864 9741 4928
rect 9805 4864 9821 4928
rect 9885 4864 9901 4928
rect 9965 4864 9973 4928
rect 9653 4863 9973 4864
rect 3121 4384 3441 4385
rect 3121 4320 3129 4384
rect 3193 4320 3209 4384
rect 3273 4320 3289 4384
rect 3353 4320 3369 4384
rect 3433 4320 3441 4384
rect 3121 4319 3441 4320
rect 7476 4384 7796 4385
rect 7476 4320 7484 4384
rect 7548 4320 7564 4384
rect 7628 4320 7644 4384
rect 7708 4320 7724 4384
rect 7788 4320 7796 4384
rect 7476 4319 7796 4320
rect 11830 4384 12150 4385
rect 11830 4320 11838 4384
rect 11902 4320 11918 4384
rect 11982 4320 11998 4384
rect 12062 4320 12078 4384
rect 12142 4320 12150 4384
rect 11830 4319 12150 4320
rect 5298 3840 5618 3841
rect 5298 3776 5306 3840
rect 5370 3776 5386 3840
rect 5450 3776 5466 3840
rect 5530 3776 5546 3840
rect 5610 3776 5618 3840
rect 5298 3775 5618 3776
rect 9653 3840 9973 3841
rect 9653 3776 9661 3840
rect 9725 3776 9741 3840
rect 9805 3776 9821 3840
rect 9885 3776 9901 3840
rect 9965 3776 9973 3840
rect 9653 3775 9973 3776
rect 3121 3296 3441 3297
rect 3121 3232 3129 3296
rect 3193 3232 3209 3296
rect 3273 3232 3289 3296
rect 3353 3232 3369 3296
rect 3433 3232 3441 3296
rect 3121 3231 3441 3232
rect 7476 3296 7796 3297
rect 7476 3232 7484 3296
rect 7548 3232 7564 3296
rect 7628 3232 7644 3296
rect 7708 3232 7724 3296
rect 7788 3232 7796 3296
rect 7476 3231 7796 3232
rect 11830 3296 12150 3297
rect 11830 3232 11838 3296
rect 11902 3232 11918 3296
rect 11982 3232 11998 3296
rect 12062 3232 12078 3296
rect 12142 3232 12150 3296
rect 11830 3231 12150 3232
rect 5298 2752 5618 2753
rect 5298 2688 5306 2752
rect 5370 2688 5386 2752
rect 5450 2688 5466 2752
rect 5530 2688 5546 2752
rect 5610 2688 5618 2752
rect 5298 2687 5618 2688
rect 9653 2752 9973 2753
rect 9653 2688 9661 2752
rect 9725 2688 9741 2752
rect 9805 2688 9821 2752
rect 9885 2688 9901 2752
rect 9965 2688 9973 2752
rect 9653 2687 9973 2688
rect 3121 2208 3441 2209
rect 3121 2144 3129 2208
rect 3193 2144 3209 2208
rect 3273 2144 3289 2208
rect 3353 2144 3369 2208
rect 3433 2144 3441 2208
rect 3121 2143 3441 2144
rect 7476 2208 7796 2209
rect 7476 2144 7484 2208
rect 7548 2144 7564 2208
rect 7628 2144 7644 2208
rect 7708 2144 7724 2208
rect 7788 2144 7796 2208
rect 7476 2143 7796 2144
rect 11830 2208 12150 2209
rect 11830 2144 11838 2208
rect 11902 2144 11918 2208
rect 11982 2144 11998 2208
rect 12062 2144 12078 2208
rect 12142 2144 12150 2208
rect 11830 2143 12150 2144
rect 13445 778 13511 781
rect 14491 778 15291 808
rect 13445 776 15291 778
rect 13445 720 13450 776
rect 13506 720 15291 776
rect 13445 718 15291 720
rect 13445 715 13511 718
rect 14491 688 15291 718
<< via3 >>
rect 3129 15260 3193 15264
rect 3129 15204 3133 15260
rect 3133 15204 3189 15260
rect 3189 15204 3193 15260
rect 3129 15200 3193 15204
rect 3209 15260 3273 15264
rect 3209 15204 3213 15260
rect 3213 15204 3269 15260
rect 3269 15204 3273 15260
rect 3209 15200 3273 15204
rect 3289 15260 3353 15264
rect 3289 15204 3293 15260
rect 3293 15204 3349 15260
rect 3349 15204 3353 15260
rect 3289 15200 3353 15204
rect 3369 15260 3433 15264
rect 3369 15204 3373 15260
rect 3373 15204 3429 15260
rect 3429 15204 3433 15260
rect 3369 15200 3433 15204
rect 7484 15260 7548 15264
rect 7484 15204 7488 15260
rect 7488 15204 7544 15260
rect 7544 15204 7548 15260
rect 7484 15200 7548 15204
rect 7564 15260 7628 15264
rect 7564 15204 7568 15260
rect 7568 15204 7624 15260
rect 7624 15204 7628 15260
rect 7564 15200 7628 15204
rect 7644 15260 7708 15264
rect 7644 15204 7648 15260
rect 7648 15204 7704 15260
rect 7704 15204 7708 15260
rect 7644 15200 7708 15204
rect 7724 15260 7788 15264
rect 7724 15204 7728 15260
rect 7728 15204 7784 15260
rect 7784 15204 7788 15260
rect 7724 15200 7788 15204
rect 11838 15260 11902 15264
rect 11838 15204 11842 15260
rect 11842 15204 11898 15260
rect 11898 15204 11902 15260
rect 11838 15200 11902 15204
rect 11918 15260 11982 15264
rect 11918 15204 11922 15260
rect 11922 15204 11978 15260
rect 11978 15204 11982 15260
rect 11918 15200 11982 15204
rect 11998 15260 12062 15264
rect 11998 15204 12002 15260
rect 12002 15204 12058 15260
rect 12058 15204 12062 15260
rect 11998 15200 12062 15204
rect 12078 15260 12142 15264
rect 12078 15204 12082 15260
rect 12082 15204 12138 15260
rect 12138 15204 12142 15260
rect 12078 15200 12142 15204
rect 5306 14716 5370 14720
rect 5306 14660 5310 14716
rect 5310 14660 5366 14716
rect 5366 14660 5370 14716
rect 5306 14656 5370 14660
rect 5386 14716 5450 14720
rect 5386 14660 5390 14716
rect 5390 14660 5446 14716
rect 5446 14660 5450 14716
rect 5386 14656 5450 14660
rect 5466 14716 5530 14720
rect 5466 14660 5470 14716
rect 5470 14660 5526 14716
rect 5526 14660 5530 14716
rect 5466 14656 5530 14660
rect 5546 14716 5610 14720
rect 5546 14660 5550 14716
rect 5550 14660 5606 14716
rect 5606 14660 5610 14716
rect 5546 14656 5610 14660
rect 9661 14716 9725 14720
rect 9661 14660 9665 14716
rect 9665 14660 9721 14716
rect 9721 14660 9725 14716
rect 9661 14656 9725 14660
rect 9741 14716 9805 14720
rect 9741 14660 9745 14716
rect 9745 14660 9801 14716
rect 9801 14660 9805 14716
rect 9741 14656 9805 14660
rect 9821 14716 9885 14720
rect 9821 14660 9825 14716
rect 9825 14660 9881 14716
rect 9881 14660 9885 14716
rect 9821 14656 9885 14660
rect 9901 14716 9965 14720
rect 9901 14660 9905 14716
rect 9905 14660 9961 14716
rect 9961 14660 9965 14716
rect 9901 14656 9965 14660
rect 3129 14172 3193 14176
rect 3129 14116 3133 14172
rect 3133 14116 3189 14172
rect 3189 14116 3193 14172
rect 3129 14112 3193 14116
rect 3209 14172 3273 14176
rect 3209 14116 3213 14172
rect 3213 14116 3269 14172
rect 3269 14116 3273 14172
rect 3209 14112 3273 14116
rect 3289 14172 3353 14176
rect 3289 14116 3293 14172
rect 3293 14116 3349 14172
rect 3349 14116 3353 14172
rect 3289 14112 3353 14116
rect 3369 14172 3433 14176
rect 3369 14116 3373 14172
rect 3373 14116 3429 14172
rect 3429 14116 3433 14172
rect 3369 14112 3433 14116
rect 7484 14172 7548 14176
rect 7484 14116 7488 14172
rect 7488 14116 7544 14172
rect 7544 14116 7548 14172
rect 7484 14112 7548 14116
rect 7564 14172 7628 14176
rect 7564 14116 7568 14172
rect 7568 14116 7624 14172
rect 7624 14116 7628 14172
rect 7564 14112 7628 14116
rect 7644 14172 7708 14176
rect 7644 14116 7648 14172
rect 7648 14116 7704 14172
rect 7704 14116 7708 14172
rect 7644 14112 7708 14116
rect 7724 14172 7788 14176
rect 7724 14116 7728 14172
rect 7728 14116 7784 14172
rect 7784 14116 7788 14172
rect 7724 14112 7788 14116
rect 11838 14172 11902 14176
rect 11838 14116 11842 14172
rect 11842 14116 11898 14172
rect 11898 14116 11902 14172
rect 11838 14112 11902 14116
rect 11918 14172 11982 14176
rect 11918 14116 11922 14172
rect 11922 14116 11978 14172
rect 11978 14116 11982 14172
rect 11918 14112 11982 14116
rect 11998 14172 12062 14176
rect 11998 14116 12002 14172
rect 12002 14116 12058 14172
rect 12058 14116 12062 14172
rect 11998 14112 12062 14116
rect 12078 14172 12142 14176
rect 12078 14116 12082 14172
rect 12082 14116 12138 14172
rect 12138 14116 12142 14172
rect 12078 14112 12142 14116
rect 5306 13628 5370 13632
rect 5306 13572 5310 13628
rect 5310 13572 5366 13628
rect 5366 13572 5370 13628
rect 5306 13568 5370 13572
rect 5386 13628 5450 13632
rect 5386 13572 5390 13628
rect 5390 13572 5446 13628
rect 5446 13572 5450 13628
rect 5386 13568 5450 13572
rect 5466 13628 5530 13632
rect 5466 13572 5470 13628
rect 5470 13572 5526 13628
rect 5526 13572 5530 13628
rect 5466 13568 5530 13572
rect 5546 13628 5610 13632
rect 5546 13572 5550 13628
rect 5550 13572 5606 13628
rect 5606 13572 5610 13628
rect 5546 13568 5610 13572
rect 9661 13628 9725 13632
rect 9661 13572 9665 13628
rect 9665 13572 9721 13628
rect 9721 13572 9725 13628
rect 9661 13568 9725 13572
rect 9741 13628 9805 13632
rect 9741 13572 9745 13628
rect 9745 13572 9801 13628
rect 9801 13572 9805 13628
rect 9741 13568 9805 13572
rect 9821 13628 9885 13632
rect 9821 13572 9825 13628
rect 9825 13572 9881 13628
rect 9881 13572 9885 13628
rect 9821 13568 9885 13572
rect 9901 13628 9965 13632
rect 9901 13572 9905 13628
rect 9905 13572 9961 13628
rect 9961 13572 9965 13628
rect 9901 13568 9965 13572
rect 3129 13084 3193 13088
rect 3129 13028 3133 13084
rect 3133 13028 3189 13084
rect 3189 13028 3193 13084
rect 3129 13024 3193 13028
rect 3209 13084 3273 13088
rect 3209 13028 3213 13084
rect 3213 13028 3269 13084
rect 3269 13028 3273 13084
rect 3209 13024 3273 13028
rect 3289 13084 3353 13088
rect 3289 13028 3293 13084
rect 3293 13028 3349 13084
rect 3349 13028 3353 13084
rect 3289 13024 3353 13028
rect 3369 13084 3433 13088
rect 3369 13028 3373 13084
rect 3373 13028 3429 13084
rect 3429 13028 3433 13084
rect 3369 13024 3433 13028
rect 7484 13084 7548 13088
rect 7484 13028 7488 13084
rect 7488 13028 7544 13084
rect 7544 13028 7548 13084
rect 7484 13024 7548 13028
rect 7564 13084 7628 13088
rect 7564 13028 7568 13084
rect 7568 13028 7624 13084
rect 7624 13028 7628 13084
rect 7564 13024 7628 13028
rect 7644 13084 7708 13088
rect 7644 13028 7648 13084
rect 7648 13028 7704 13084
rect 7704 13028 7708 13084
rect 7644 13024 7708 13028
rect 7724 13084 7788 13088
rect 7724 13028 7728 13084
rect 7728 13028 7784 13084
rect 7784 13028 7788 13084
rect 7724 13024 7788 13028
rect 11838 13084 11902 13088
rect 11838 13028 11842 13084
rect 11842 13028 11898 13084
rect 11898 13028 11902 13084
rect 11838 13024 11902 13028
rect 11918 13084 11982 13088
rect 11918 13028 11922 13084
rect 11922 13028 11978 13084
rect 11978 13028 11982 13084
rect 11918 13024 11982 13028
rect 11998 13084 12062 13088
rect 11998 13028 12002 13084
rect 12002 13028 12058 13084
rect 12058 13028 12062 13084
rect 11998 13024 12062 13028
rect 12078 13084 12142 13088
rect 12078 13028 12082 13084
rect 12082 13028 12138 13084
rect 12138 13028 12142 13084
rect 12078 13024 12142 13028
rect 5306 12540 5370 12544
rect 5306 12484 5310 12540
rect 5310 12484 5366 12540
rect 5366 12484 5370 12540
rect 5306 12480 5370 12484
rect 5386 12540 5450 12544
rect 5386 12484 5390 12540
rect 5390 12484 5446 12540
rect 5446 12484 5450 12540
rect 5386 12480 5450 12484
rect 5466 12540 5530 12544
rect 5466 12484 5470 12540
rect 5470 12484 5526 12540
rect 5526 12484 5530 12540
rect 5466 12480 5530 12484
rect 5546 12540 5610 12544
rect 5546 12484 5550 12540
rect 5550 12484 5606 12540
rect 5606 12484 5610 12540
rect 5546 12480 5610 12484
rect 9661 12540 9725 12544
rect 9661 12484 9665 12540
rect 9665 12484 9721 12540
rect 9721 12484 9725 12540
rect 9661 12480 9725 12484
rect 9741 12540 9805 12544
rect 9741 12484 9745 12540
rect 9745 12484 9801 12540
rect 9801 12484 9805 12540
rect 9741 12480 9805 12484
rect 9821 12540 9885 12544
rect 9821 12484 9825 12540
rect 9825 12484 9881 12540
rect 9881 12484 9885 12540
rect 9821 12480 9885 12484
rect 9901 12540 9965 12544
rect 9901 12484 9905 12540
rect 9905 12484 9961 12540
rect 9961 12484 9965 12540
rect 9901 12480 9965 12484
rect 3129 11996 3193 12000
rect 3129 11940 3133 11996
rect 3133 11940 3189 11996
rect 3189 11940 3193 11996
rect 3129 11936 3193 11940
rect 3209 11996 3273 12000
rect 3209 11940 3213 11996
rect 3213 11940 3269 11996
rect 3269 11940 3273 11996
rect 3209 11936 3273 11940
rect 3289 11996 3353 12000
rect 3289 11940 3293 11996
rect 3293 11940 3349 11996
rect 3349 11940 3353 11996
rect 3289 11936 3353 11940
rect 3369 11996 3433 12000
rect 3369 11940 3373 11996
rect 3373 11940 3429 11996
rect 3429 11940 3433 11996
rect 3369 11936 3433 11940
rect 7484 11996 7548 12000
rect 7484 11940 7488 11996
rect 7488 11940 7544 11996
rect 7544 11940 7548 11996
rect 7484 11936 7548 11940
rect 7564 11996 7628 12000
rect 7564 11940 7568 11996
rect 7568 11940 7624 11996
rect 7624 11940 7628 11996
rect 7564 11936 7628 11940
rect 7644 11996 7708 12000
rect 7644 11940 7648 11996
rect 7648 11940 7704 11996
rect 7704 11940 7708 11996
rect 7644 11936 7708 11940
rect 7724 11996 7788 12000
rect 7724 11940 7728 11996
rect 7728 11940 7784 11996
rect 7784 11940 7788 11996
rect 7724 11936 7788 11940
rect 11838 11996 11902 12000
rect 11838 11940 11842 11996
rect 11842 11940 11898 11996
rect 11898 11940 11902 11996
rect 11838 11936 11902 11940
rect 11918 11996 11982 12000
rect 11918 11940 11922 11996
rect 11922 11940 11978 11996
rect 11978 11940 11982 11996
rect 11918 11936 11982 11940
rect 11998 11996 12062 12000
rect 11998 11940 12002 11996
rect 12002 11940 12058 11996
rect 12058 11940 12062 11996
rect 11998 11936 12062 11940
rect 12078 11996 12142 12000
rect 12078 11940 12082 11996
rect 12082 11940 12138 11996
rect 12138 11940 12142 11996
rect 12078 11936 12142 11940
rect 5306 11452 5370 11456
rect 5306 11396 5310 11452
rect 5310 11396 5366 11452
rect 5366 11396 5370 11452
rect 5306 11392 5370 11396
rect 5386 11452 5450 11456
rect 5386 11396 5390 11452
rect 5390 11396 5446 11452
rect 5446 11396 5450 11452
rect 5386 11392 5450 11396
rect 5466 11452 5530 11456
rect 5466 11396 5470 11452
rect 5470 11396 5526 11452
rect 5526 11396 5530 11452
rect 5466 11392 5530 11396
rect 5546 11452 5610 11456
rect 5546 11396 5550 11452
rect 5550 11396 5606 11452
rect 5606 11396 5610 11452
rect 5546 11392 5610 11396
rect 9661 11452 9725 11456
rect 9661 11396 9665 11452
rect 9665 11396 9721 11452
rect 9721 11396 9725 11452
rect 9661 11392 9725 11396
rect 9741 11452 9805 11456
rect 9741 11396 9745 11452
rect 9745 11396 9801 11452
rect 9801 11396 9805 11452
rect 9741 11392 9805 11396
rect 9821 11452 9885 11456
rect 9821 11396 9825 11452
rect 9825 11396 9881 11452
rect 9881 11396 9885 11452
rect 9821 11392 9885 11396
rect 9901 11452 9965 11456
rect 9901 11396 9905 11452
rect 9905 11396 9961 11452
rect 9961 11396 9965 11452
rect 9901 11392 9965 11396
rect 3129 10908 3193 10912
rect 3129 10852 3133 10908
rect 3133 10852 3189 10908
rect 3189 10852 3193 10908
rect 3129 10848 3193 10852
rect 3209 10908 3273 10912
rect 3209 10852 3213 10908
rect 3213 10852 3269 10908
rect 3269 10852 3273 10908
rect 3209 10848 3273 10852
rect 3289 10908 3353 10912
rect 3289 10852 3293 10908
rect 3293 10852 3349 10908
rect 3349 10852 3353 10908
rect 3289 10848 3353 10852
rect 3369 10908 3433 10912
rect 3369 10852 3373 10908
rect 3373 10852 3429 10908
rect 3429 10852 3433 10908
rect 3369 10848 3433 10852
rect 7484 10908 7548 10912
rect 7484 10852 7488 10908
rect 7488 10852 7544 10908
rect 7544 10852 7548 10908
rect 7484 10848 7548 10852
rect 7564 10908 7628 10912
rect 7564 10852 7568 10908
rect 7568 10852 7624 10908
rect 7624 10852 7628 10908
rect 7564 10848 7628 10852
rect 7644 10908 7708 10912
rect 7644 10852 7648 10908
rect 7648 10852 7704 10908
rect 7704 10852 7708 10908
rect 7644 10848 7708 10852
rect 7724 10908 7788 10912
rect 7724 10852 7728 10908
rect 7728 10852 7784 10908
rect 7784 10852 7788 10908
rect 7724 10848 7788 10852
rect 11838 10908 11902 10912
rect 11838 10852 11842 10908
rect 11842 10852 11898 10908
rect 11898 10852 11902 10908
rect 11838 10848 11902 10852
rect 11918 10908 11982 10912
rect 11918 10852 11922 10908
rect 11922 10852 11978 10908
rect 11978 10852 11982 10908
rect 11918 10848 11982 10852
rect 11998 10908 12062 10912
rect 11998 10852 12002 10908
rect 12002 10852 12058 10908
rect 12058 10852 12062 10908
rect 11998 10848 12062 10852
rect 12078 10908 12142 10912
rect 12078 10852 12082 10908
rect 12082 10852 12138 10908
rect 12138 10852 12142 10908
rect 12078 10848 12142 10852
rect 5306 10364 5370 10368
rect 5306 10308 5310 10364
rect 5310 10308 5366 10364
rect 5366 10308 5370 10364
rect 5306 10304 5370 10308
rect 5386 10364 5450 10368
rect 5386 10308 5390 10364
rect 5390 10308 5446 10364
rect 5446 10308 5450 10364
rect 5386 10304 5450 10308
rect 5466 10364 5530 10368
rect 5466 10308 5470 10364
rect 5470 10308 5526 10364
rect 5526 10308 5530 10364
rect 5466 10304 5530 10308
rect 5546 10364 5610 10368
rect 5546 10308 5550 10364
rect 5550 10308 5606 10364
rect 5606 10308 5610 10364
rect 5546 10304 5610 10308
rect 9661 10364 9725 10368
rect 9661 10308 9665 10364
rect 9665 10308 9721 10364
rect 9721 10308 9725 10364
rect 9661 10304 9725 10308
rect 9741 10364 9805 10368
rect 9741 10308 9745 10364
rect 9745 10308 9801 10364
rect 9801 10308 9805 10364
rect 9741 10304 9805 10308
rect 9821 10364 9885 10368
rect 9821 10308 9825 10364
rect 9825 10308 9881 10364
rect 9881 10308 9885 10364
rect 9821 10304 9885 10308
rect 9901 10364 9965 10368
rect 9901 10308 9905 10364
rect 9905 10308 9961 10364
rect 9961 10308 9965 10364
rect 9901 10304 9965 10308
rect 3129 9820 3193 9824
rect 3129 9764 3133 9820
rect 3133 9764 3189 9820
rect 3189 9764 3193 9820
rect 3129 9760 3193 9764
rect 3209 9820 3273 9824
rect 3209 9764 3213 9820
rect 3213 9764 3269 9820
rect 3269 9764 3273 9820
rect 3209 9760 3273 9764
rect 3289 9820 3353 9824
rect 3289 9764 3293 9820
rect 3293 9764 3349 9820
rect 3349 9764 3353 9820
rect 3289 9760 3353 9764
rect 3369 9820 3433 9824
rect 3369 9764 3373 9820
rect 3373 9764 3429 9820
rect 3429 9764 3433 9820
rect 3369 9760 3433 9764
rect 7484 9820 7548 9824
rect 7484 9764 7488 9820
rect 7488 9764 7544 9820
rect 7544 9764 7548 9820
rect 7484 9760 7548 9764
rect 7564 9820 7628 9824
rect 7564 9764 7568 9820
rect 7568 9764 7624 9820
rect 7624 9764 7628 9820
rect 7564 9760 7628 9764
rect 7644 9820 7708 9824
rect 7644 9764 7648 9820
rect 7648 9764 7704 9820
rect 7704 9764 7708 9820
rect 7644 9760 7708 9764
rect 7724 9820 7788 9824
rect 7724 9764 7728 9820
rect 7728 9764 7784 9820
rect 7784 9764 7788 9820
rect 7724 9760 7788 9764
rect 11838 9820 11902 9824
rect 11838 9764 11842 9820
rect 11842 9764 11898 9820
rect 11898 9764 11902 9820
rect 11838 9760 11902 9764
rect 11918 9820 11982 9824
rect 11918 9764 11922 9820
rect 11922 9764 11978 9820
rect 11978 9764 11982 9820
rect 11918 9760 11982 9764
rect 11998 9820 12062 9824
rect 11998 9764 12002 9820
rect 12002 9764 12058 9820
rect 12058 9764 12062 9820
rect 11998 9760 12062 9764
rect 12078 9820 12142 9824
rect 12078 9764 12082 9820
rect 12082 9764 12138 9820
rect 12138 9764 12142 9820
rect 12078 9760 12142 9764
rect 5306 9276 5370 9280
rect 5306 9220 5310 9276
rect 5310 9220 5366 9276
rect 5366 9220 5370 9276
rect 5306 9216 5370 9220
rect 5386 9276 5450 9280
rect 5386 9220 5390 9276
rect 5390 9220 5446 9276
rect 5446 9220 5450 9276
rect 5386 9216 5450 9220
rect 5466 9276 5530 9280
rect 5466 9220 5470 9276
rect 5470 9220 5526 9276
rect 5526 9220 5530 9276
rect 5466 9216 5530 9220
rect 5546 9276 5610 9280
rect 5546 9220 5550 9276
rect 5550 9220 5606 9276
rect 5606 9220 5610 9276
rect 5546 9216 5610 9220
rect 9661 9276 9725 9280
rect 9661 9220 9665 9276
rect 9665 9220 9721 9276
rect 9721 9220 9725 9276
rect 9661 9216 9725 9220
rect 9741 9276 9805 9280
rect 9741 9220 9745 9276
rect 9745 9220 9801 9276
rect 9801 9220 9805 9276
rect 9741 9216 9805 9220
rect 9821 9276 9885 9280
rect 9821 9220 9825 9276
rect 9825 9220 9881 9276
rect 9881 9220 9885 9276
rect 9821 9216 9885 9220
rect 9901 9276 9965 9280
rect 9901 9220 9905 9276
rect 9905 9220 9961 9276
rect 9961 9220 9965 9276
rect 9901 9216 9965 9220
rect 3129 8732 3193 8736
rect 3129 8676 3133 8732
rect 3133 8676 3189 8732
rect 3189 8676 3193 8732
rect 3129 8672 3193 8676
rect 3209 8732 3273 8736
rect 3209 8676 3213 8732
rect 3213 8676 3269 8732
rect 3269 8676 3273 8732
rect 3209 8672 3273 8676
rect 3289 8732 3353 8736
rect 3289 8676 3293 8732
rect 3293 8676 3349 8732
rect 3349 8676 3353 8732
rect 3289 8672 3353 8676
rect 3369 8732 3433 8736
rect 3369 8676 3373 8732
rect 3373 8676 3429 8732
rect 3429 8676 3433 8732
rect 3369 8672 3433 8676
rect 7484 8732 7548 8736
rect 7484 8676 7488 8732
rect 7488 8676 7544 8732
rect 7544 8676 7548 8732
rect 7484 8672 7548 8676
rect 7564 8732 7628 8736
rect 7564 8676 7568 8732
rect 7568 8676 7624 8732
rect 7624 8676 7628 8732
rect 7564 8672 7628 8676
rect 7644 8732 7708 8736
rect 7644 8676 7648 8732
rect 7648 8676 7704 8732
rect 7704 8676 7708 8732
rect 7644 8672 7708 8676
rect 7724 8732 7788 8736
rect 7724 8676 7728 8732
rect 7728 8676 7784 8732
rect 7784 8676 7788 8732
rect 7724 8672 7788 8676
rect 11838 8732 11902 8736
rect 11838 8676 11842 8732
rect 11842 8676 11898 8732
rect 11898 8676 11902 8732
rect 11838 8672 11902 8676
rect 11918 8732 11982 8736
rect 11918 8676 11922 8732
rect 11922 8676 11978 8732
rect 11978 8676 11982 8732
rect 11918 8672 11982 8676
rect 11998 8732 12062 8736
rect 11998 8676 12002 8732
rect 12002 8676 12058 8732
rect 12058 8676 12062 8732
rect 11998 8672 12062 8676
rect 12078 8732 12142 8736
rect 12078 8676 12082 8732
rect 12082 8676 12138 8732
rect 12138 8676 12142 8732
rect 12078 8672 12142 8676
rect 5306 8188 5370 8192
rect 5306 8132 5310 8188
rect 5310 8132 5366 8188
rect 5366 8132 5370 8188
rect 5306 8128 5370 8132
rect 5386 8188 5450 8192
rect 5386 8132 5390 8188
rect 5390 8132 5446 8188
rect 5446 8132 5450 8188
rect 5386 8128 5450 8132
rect 5466 8188 5530 8192
rect 5466 8132 5470 8188
rect 5470 8132 5526 8188
rect 5526 8132 5530 8188
rect 5466 8128 5530 8132
rect 5546 8188 5610 8192
rect 5546 8132 5550 8188
rect 5550 8132 5606 8188
rect 5606 8132 5610 8188
rect 5546 8128 5610 8132
rect 9661 8188 9725 8192
rect 9661 8132 9665 8188
rect 9665 8132 9721 8188
rect 9721 8132 9725 8188
rect 9661 8128 9725 8132
rect 9741 8188 9805 8192
rect 9741 8132 9745 8188
rect 9745 8132 9801 8188
rect 9801 8132 9805 8188
rect 9741 8128 9805 8132
rect 9821 8188 9885 8192
rect 9821 8132 9825 8188
rect 9825 8132 9881 8188
rect 9881 8132 9885 8188
rect 9821 8128 9885 8132
rect 9901 8188 9965 8192
rect 9901 8132 9905 8188
rect 9905 8132 9961 8188
rect 9961 8132 9965 8188
rect 9901 8128 9965 8132
rect 3129 7644 3193 7648
rect 3129 7588 3133 7644
rect 3133 7588 3189 7644
rect 3189 7588 3193 7644
rect 3129 7584 3193 7588
rect 3209 7644 3273 7648
rect 3209 7588 3213 7644
rect 3213 7588 3269 7644
rect 3269 7588 3273 7644
rect 3209 7584 3273 7588
rect 3289 7644 3353 7648
rect 3289 7588 3293 7644
rect 3293 7588 3349 7644
rect 3349 7588 3353 7644
rect 3289 7584 3353 7588
rect 3369 7644 3433 7648
rect 3369 7588 3373 7644
rect 3373 7588 3429 7644
rect 3429 7588 3433 7644
rect 3369 7584 3433 7588
rect 7484 7644 7548 7648
rect 7484 7588 7488 7644
rect 7488 7588 7544 7644
rect 7544 7588 7548 7644
rect 7484 7584 7548 7588
rect 7564 7644 7628 7648
rect 7564 7588 7568 7644
rect 7568 7588 7624 7644
rect 7624 7588 7628 7644
rect 7564 7584 7628 7588
rect 7644 7644 7708 7648
rect 7644 7588 7648 7644
rect 7648 7588 7704 7644
rect 7704 7588 7708 7644
rect 7644 7584 7708 7588
rect 7724 7644 7788 7648
rect 7724 7588 7728 7644
rect 7728 7588 7784 7644
rect 7784 7588 7788 7644
rect 7724 7584 7788 7588
rect 11838 7644 11902 7648
rect 11838 7588 11842 7644
rect 11842 7588 11898 7644
rect 11898 7588 11902 7644
rect 11838 7584 11902 7588
rect 11918 7644 11982 7648
rect 11918 7588 11922 7644
rect 11922 7588 11978 7644
rect 11978 7588 11982 7644
rect 11918 7584 11982 7588
rect 11998 7644 12062 7648
rect 11998 7588 12002 7644
rect 12002 7588 12058 7644
rect 12058 7588 12062 7644
rect 11998 7584 12062 7588
rect 12078 7644 12142 7648
rect 12078 7588 12082 7644
rect 12082 7588 12138 7644
rect 12138 7588 12142 7644
rect 12078 7584 12142 7588
rect 5306 7100 5370 7104
rect 5306 7044 5310 7100
rect 5310 7044 5366 7100
rect 5366 7044 5370 7100
rect 5306 7040 5370 7044
rect 5386 7100 5450 7104
rect 5386 7044 5390 7100
rect 5390 7044 5446 7100
rect 5446 7044 5450 7100
rect 5386 7040 5450 7044
rect 5466 7100 5530 7104
rect 5466 7044 5470 7100
rect 5470 7044 5526 7100
rect 5526 7044 5530 7100
rect 5466 7040 5530 7044
rect 5546 7100 5610 7104
rect 5546 7044 5550 7100
rect 5550 7044 5606 7100
rect 5606 7044 5610 7100
rect 5546 7040 5610 7044
rect 9661 7100 9725 7104
rect 9661 7044 9665 7100
rect 9665 7044 9721 7100
rect 9721 7044 9725 7100
rect 9661 7040 9725 7044
rect 9741 7100 9805 7104
rect 9741 7044 9745 7100
rect 9745 7044 9801 7100
rect 9801 7044 9805 7100
rect 9741 7040 9805 7044
rect 9821 7100 9885 7104
rect 9821 7044 9825 7100
rect 9825 7044 9881 7100
rect 9881 7044 9885 7100
rect 9821 7040 9885 7044
rect 9901 7100 9965 7104
rect 9901 7044 9905 7100
rect 9905 7044 9961 7100
rect 9961 7044 9965 7100
rect 9901 7040 9965 7044
rect 3129 6556 3193 6560
rect 3129 6500 3133 6556
rect 3133 6500 3189 6556
rect 3189 6500 3193 6556
rect 3129 6496 3193 6500
rect 3209 6556 3273 6560
rect 3209 6500 3213 6556
rect 3213 6500 3269 6556
rect 3269 6500 3273 6556
rect 3209 6496 3273 6500
rect 3289 6556 3353 6560
rect 3289 6500 3293 6556
rect 3293 6500 3349 6556
rect 3349 6500 3353 6556
rect 3289 6496 3353 6500
rect 3369 6556 3433 6560
rect 3369 6500 3373 6556
rect 3373 6500 3429 6556
rect 3429 6500 3433 6556
rect 3369 6496 3433 6500
rect 7484 6556 7548 6560
rect 7484 6500 7488 6556
rect 7488 6500 7544 6556
rect 7544 6500 7548 6556
rect 7484 6496 7548 6500
rect 7564 6556 7628 6560
rect 7564 6500 7568 6556
rect 7568 6500 7624 6556
rect 7624 6500 7628 6556
rect 7564 6496 7628 6500
rect 7644 6556 7708 6560
rect 7644 6500 7648 6556
rect 7648 6500 7704 6556
rect 7704 6500 7708 6556
rect 7644 6496 7708 6500
rect 7724 6556 7788 6560
rect 7724 6500 7728 6556
rect 7728 6500 7784 6556
rect 7784 6500 7788 6556
rect 7724 6496 7788 6500
rect 11838 6556 11902 6560
rect 11838 6500 11842 6556
rect 11842 6500 11898 6556
rect 11898 6500 11902 6556
rect 11838 6496 11902 6500
rect 11918 6556 11982 6560
rect 11918 6500 11922 6556
rect 11922 6500 11978 6556
rect 11978 6500 11982 6556
rect 11918 6496 11982 6500
rect 11998 6556 12062 6560
rect 11998 6500 12002 6556
rect 12002 6500 12058 6556
rect 12058 6500 12062 6556
rect 11998 6496 12062 6500
rect 12078 6556 12142 6560
rect 12078 6500 12082 6556
rect 12082 6500 12138 6556
rect 12138 6500 12142 6556
rect 12078 6496 12142 6500
rect 5306 6012 5370 6016
rect 5306 5956 5310 6012
rect 5310 5956 5366 6012
rect 5366 5956 5370 6012
rect 5306 5952 5370 5956
rect 5386 6012 5450 6016
rect 5386 5956 5390 6012
rect 5390 5956 5446 6012
rect 5446 5956 5450 6012
rect 5386 5952 5450 5956
rect 5466 6012 5530 6016
rect 5466 5956 5470 6012
rect 5470 5956 5526 6012
rect 5526 5956 5530 6012
rect 5466 5952 5530 5956
rect 5546 6012 5610 6016
rect 5546 5956 5550 6012
rect 5550 5956 5606 6012
rect 5606 5956 5610 6012
rect 5546 5952 5610 5956
rect 9661 6012 9725 6016
rect 9661 5956 9665 6012
rect 9665 5956 9721 6012
rect 9721 5956 9725 6012
rect 9661 5952 9725 5956
rect 9741 6012 9805 6016
rect 9741 5956 9745 6012
rect 9745 5956 9801 6012
rect 9801 5956 9805 6012
rect 9741 5952 9805 5956
rect 9821 6012 9885 6016
rect 9821 5956 9825 6012
rect 9825 5956 9881 6012
rect 9881 5956 9885 6012
rect 9821 5952 9885 5956
rect 9901 6012 9965 6016
rect 9901 5956 9905 6012
rect 9905 5956 9961 6012
rect 9961 5956 9965 6012
rect 9901 5952 9965 5956
rect 3129 5468 3193 5472
rect 3129 5412 3133 5468
rect 3133 5412 3189 5468
rect 3189 5412 3193 5468
rect 3129 5408 3193 5412
rect 3209 5468 3273 5472
rect 3209 5412 3213 5468
rect 3213 5412 3269 5468
rect 3269 5412 3273 5468
rect 3209 5408 3273 5412
rect 3289 5468 3353 5472
rect 3289 5412 3293 5468
rect 3293 5412 3349 5468
rect 3349 5412 3353 5468
rect 3289 5408 3353 5412
rect 3369 5468 3433 5472
rect 3369 5412 3373 5468
rect 3373 5412 3429 5468
rect 3429 5412 3433 5468
rect 3369 5408 3433 5412
rect 7484 5468 7548 5472
rect 7484 5412 7488 5468
rect 7488 5412 7544 5468
rect 7544 5412 7548 5468
rect 7484 5408 7548 5412
rect 7564 5468 7628 5472
rect 7564 5412 7568 5468
rect 7568 5412 7624 5468
rect 7624 5412 7628 5468
rect 7564 5408 7628 5412
rect 7644 5468 7708 5472
rect 7644 5412 7648 5468
rect 7648 5412 7704 5468
rect 7704 5412 7708 5468
rect 7644 5408 7708 5412
rect 7724 5468 7788 5472
rect 7724 5412 7728 5468
rect 7728 5412 7784 5468
rect 7784 5412 7788 5468
rect 7724 5408 7788 5412
rect 11838 5468 11902 5472
rect 11838 5412 11842 5468
rect 11842 5412 11898 5468
rect 11898 5412 11902 5468
rect 11838 5408 11902 5412
rect 11918 5468 11982 5472
rect 11918 5412 11922 5468
rect 11922 5412 11978 5468
rect 11978 5412 11982 5468
rect 11918 5408 11982 5412
rect 11998 5468 12062 5472
rect 11998 5412 12002 5468
rect 12002 5412 12058 5468
rect 12058 5412 12062 5468
rect 11998 5408 12062 5412
rect 12078 5468 12142 5472
rect 12078 5412 12082 5468
rect 12082 5412 12138 5468
rect 12138 5412 12142 5468
rect 12078 5408 12142 5412
rect 5306 4924 5370 4928
rect 5306 4868 5310 4924
rect 5310 4868 5366 4924
rect 5366 4868 5370 4924
rect 5306 4864 5370 4868
rect 5386 4924 5450 4928
rect 5386 4868 5390 4924
rect 5390 4868 5446 4924
rect 5446 4868 5450 4924
rect 5386 4864 5450 4868
rect 5466 4924 5530 4928
rect 5466 4868 5470 4924
rect 5470 4868 5526 4924
rect 5526 4868 5530 4924
rect 5466 4864 5530 4868
rect 5546 4924 5610 4928
rect 5546 4868 5550 4924
rect 5550 4868 5606 4924
rect 5606 4868 5610 4924
rect 5546 4864 5610 4868
rect 9661 4924 9725 4928
rect 9661 4868 9665 4924
rect 9665 4868 9721 4924
rect 9721 4868 9725 4924
rect 9661 4864 9725 4868
rect 9741 4924 9805 4928
rect 9741 4868 9745 4924
rect 9745 4868 9801 4924
rect 9801 4868 9805 4924
rect 9741 4864 9805 4868
rect 9821 4924 9885 4928
rect 9821 4868 9825 4924
rect 9825 4868 9881 4924
rect 9881 4868 9885 4924
rect 9821 4864 9885 4868
rect 9901 4924 9965 4928
rect 9901 4868 9905 4924
rect 9905 4868 9961 4924
rect 9961 4868 9965 4924
rect 9901 4864 9965 4868
rect 3129 4380 3193 4384
rect 3129 4324 3133 4380
rect 3133 4324 3189 4380
rect 3189 4324 3193 4380
rect 3129 4320 3193 4324
rect 3209 4380 3273 4384
rect 3209 4324 3213 4380
rect 3213 4324 3269 4380
rect 3269 4324 3273 4380
rect 3209 4320 3273 4324
rect 3289 4380 3353 4384
rect 3289 4324 3293 4380
rect 3293 4324 3349 4380
rect 3349 4324 3353 4380
rect 3289 4320 3353 4324
rect 3369 4380 3433 4384
rect 3369 4324 3373 4380
rect 3373 4324 3429 4380
rect 3429 4324 3433 4380
rect 3369 4320 3433 4324
rect 7484 4380 7548 4384
rect 7484 4324 7488 4380
rect 7488 4324 7544 4380
rect 7544 4324 7548 4380
rect 7484 4320 7548 4324
rect 7564 4380 7628 4384
rect 7564 4324 7568 4380
rect 7568 4324 7624 4380
rect 7624 4324 7628 4380
rect 7564 4320 7628 4324
rect 7644 4380 7708 4384
rect 7644 4324 7648 4380
rect 7648 4324 7704 4380
rect 7704 4324 7708 4380
rect 7644 4320 7708 4324
rect 7724 4380 7788 4384
rect 7724 4324 7728 4380
rect 7728 4324 7784 4380
rect 7784 4324 7788 4380
rect 7724 4320 7788 4324
rect 11838 4380 11902 4384
rect 11838 4324 11842 4380
rect 11842 4324 11898 4380
rect 11898 4324 11902 4380
rect 11838 4320 11902 4324
rect 11918 4380 11982 4384
rect 11918 4324 11922 4380
rect 11922 4324 11978 4380
rect 11978 4324 11982 4380
rect 11918 4320 11982 4324
rect 11998 4380 12062 4384
rect 11998 4324 12002 4380
rect 12002 4324 12058 4380
rect 12058 4324 12062 4380
rect 11998 4320 12062 4324
rect 12078 4380 12142 4384
rect 12078 4324 12082 4380
rect 12082 4324 12138 4380
rect 12138 4324 12142 4380
rect 12078 4320 12142 4324
rect 5306 3836 5370 3840
rect 5306 3780 5310 3836
rect 5310 3780 5366 3836
rect 5366 3780 5370 3836
rect 5306 3776 5370 3780
rect 5386 3836 5450 3840
rect 5386 3780 5390 3836
rect 5390 3780 5446 3836
rect 5446 3780 5450 3836
rect 5386 3776 5450 3780
rect 5466 3836 5530 3840
rect 5466 3780 5470 3836
rect 5470 3780 5526 3836
rect 5526 3780 5530 3836
rect 5466 3776 5530 3780
rect 5546 3836 5610 3840
rect 5546 3780 5550 3836
rect 5550 3780 5606 3836
rect 5606 3780 5610 3836
rect 5546 3776 5610 3780
rect 9661 3836 9725 3840
rect 9661 3780 9665 3836
rect 9665 3780 9721 3836
rect 9721 3780 9725 3836
rect 9661 3776 9725 3780
rect 9741 3836 9805 3840
rect 9741 3780 9745 3836
rect 9745 3780 9801 3836
rect 9801 3780 9805 3836
rect 9741 3776 9805 3780
rect 9821 3836 9885 3840
rect 9821 3780 9825 3836
rect 9825 3780 9881 3836
rect 9881 3780 9885 3836
rect 9821 3776 9885 3780
rect 9901 3836 9965 3840
rect 9901 3780 9905 3836
rect 9905 3780 9961 3836
rect 9961 3780 9965 3836
rect 9901 3776 9965 3780
rect 3129 3292 3193 3296
rect 3129 3236 3133 3292
rect 3133 3236 3189 3292
rect 3189 3236 3193 3292
rect 3129 3232 3193 3236
rect 3209 3292 3273 3296
rect 3209 3236 3213 3292
rect 3213 3236 3269 3292
rect 3269 3236 3273 3292
rect 3209 3232 3273 3236
rect 3289 3292 3353 3296
rect 3289 3236 3293 3292
rect 3293 3236 3349 3292
rect 3349 3236 3353 3292
rect 3289 3232 3353 3236
rect 3369 3292 3433 3296
rect 3369 3236 3373 3292
rect 3373 3236 3429 3292
rect 3429 3236 3433 3292
rect 3369 3232 3433 3236
rect 7484 3292 7548 3296
rect 7484 3236 7488 3292
rect 7488 3236 7544 3292
rect 7544 3236 7548 3292
rect 7484 3232 7548 3236
rect 7564 3292 7628 3296
rect 7564 3236 7568 3292
rect 7568 3236 7624 3292
rect 7624 3236 7628 3292
rect 7564 3232 7628 3236
rect 7644 3292 7708 3296
rect 7644 3236 7648 3292
rect 7648 3236 7704 3292
rect 7704 3236 7708 3292
rect 7644 3232 7708 3236
rect 7724 3292 7788 3296
rect 7724 3236 7728 3292
rect 7728 3236 7784 3292
rect 7784 3236 7788 3292
rect 7724 3232 7788 3236
rect 11838 3292 11902 3296
rect 11838 3236 11842 3292
rect 11842 3236 11898 3292
rect 11898 3236 11902 3292
rect 11838 3232 11902 3236
rect 11918 3292 11982 3296
rect 11918 3236 11922 3292
rect 11922 3236 11978 3292
rect 11978 3236 11982 3292
rect 11918 3232 11982 3236
rect 11998 3292 12062 3296
rect 11998 3236 12002 3292
rect 12002 3236 12058 3292
rect 12058 3236 12062 3292
rect 11998 3232 12062 3236
rect 12078 3292 12142 3296
rect 12078 3236 12082 3292
rect 12082 3236 12138 3292
rect 12138 3236 12142 3292
rect 12078 3232 12142 3236
rect 5306 2748 5370 2752
rect 5306 2692 5310 2748
rect 5310 2692 5366 2748
rect 5366 2692 5370 2748
rect 5306 2688 5370 2692
rect 5386 2748 5450 2752
rect 5386 2692 5390 2748
rect 5390 2692 5446 2748
rect 5446 2692 5450 2748
rect 5386 2688 5450 2692
rect 5466 2748 5530 2752
rect 5466 2692 5470 2748
rect 5470 2692 5526 2748
rect 5526 2692 5530 2748
rect 5466 2688 5530 2692
rect 5546 2748 5610 2752
rect 5546 2692 5550 2748
rect 5550 2692 5606 2748
rect 5606 2692 5610 2748
rect 5546 2688 5610 2692
rect 9661 2748 9725 2752
rect 9661 2692 9665 2748
rect 9665 2692 9721 2748
rect 9721 2692 9725 2748
rect 9661 2688 9725 2692
rect 9741 2748 9805 2752
rect 9741 2692 9745 2748
rect 9745 2692 9801 2748
rect 9801 2692 9805 2748
rect 9741 2688 9805 2692
rect 9821 2748 9885 2752
rect 9821 2692 9825 2748
rect 9825 2692 9881 2748
rect 9881 2692 9885 2748
rect 9821 2688 9885 2692
rect 9901 2748 9965 2752
rect 9901 2692 9905 2748
rect 9905 2692 9961 2748
rect 9961 2692 9965 2748
rect 9901 2688 9965 2692
rect 3129 2204 3193 2208
rect 3129 2148 3133 2204
rect 3133 2148 3189 2204
rect 3189 2148 3193 2204
rect 3129 2144 3193 2148
rect 3209 2204 3273 2208
rect 3209 2148 3213 2204
rect 3213 2148 3269 2204
rect 3269 2148 3273 2204
rect 3209 2144 3273 2148
rect 3289 2204 3353 2208
rect 3289 2148 3293 2204
rect 3293 2148 3349 2204
rect 3349 2148 3353 2204
rect 3289 2144 3353 2148
rect 3369 2204 3433 2208
rect 3369 2148 3373 2204
rect 3373 2148 3429 2204
rect 3429 2148 3433 2204
rect 3369 2144 3433 2148
rect 7484 2204 7548 2208
rect 7484 2148 7488 2204
rect 7488 2148 7544 2204
rect 7544 2148 7548 2204
rect 7484 2144 7548 2148
rect 7564 2204 7628 2208
rect 7564 2148 7568 2204
rect 7568 2148 7624 2204
rect 7624 2148 7628 2204
rect 7564 2144 7628 2148
rect 7644 2204 7708 2208
rect 7644 2148 7648 2204
rect 7648 2148 7704 2204
rect 7704 2148 7708 2204
rect 7644 2144 7708 2148
rect 7724 2204 7788 2208
rect 7724 2148 7728 2204
rect 7728 2148 7784 2204
rect 7784 2148 7788 2204
rect 7724 2144 7788 2148
rect 11838 2204 11902 2208
rect 11838 2148 11842 2204
rect 11842 2148 11898 2204
rect 11898 2148 11902 2204
rect 11838 2144 11902 2148
rect 11918 2204 11982 2208
rect 11918 2148 11922 2204
rect 11922 2148 11978 2204
rect 11978 2148 11982 2204
rect 11918 2144 11982 2148
rect 11998 2204 12062 2208
rect 11998 2148 12002 2204
rect 12002 2148 12058 2204
rect 12058 2148 12062 2204
rect 11998 2144 12062 2148
rect 12078 2204 12142 2208
rect 12078 2148 12082 2204
rect 12082 2148 12138 2204
rect 12138 2148 12142 2204
rect 12078 2144 12142 2148
<< metal4 >>
rect 3121 15264 3441 15280
rect 3121 15200 3129 15264
rect 3193 15200 3209 15264
rect 3273 15200 3289 15264
rect 3353 15200 3369 15264
rect 3433 15200 3441 15264
rect 3121 14176 3441 15200
rect 3121 14112 3129 14176
rect 3193 14112 3209 14176
rect 3273 14112 3289 14176
rect 3353 14112 3369 14176
rect 3433 14112 3441 14176
rect 3121 13126 3441 14112
rect 3121 13088 3163 13126
rect 3399 13088 3441 13126
rect 3121 13024 3129 13088
rect 3433 13024 3441 13088
rect 3121 12890 3163 13024
rect 3399 12890 3441 13024
rect 3121 12000 3441 12890
rect 3121 11936 3129 12000
rect 3193 11936 3209 12000
rect 3273 11936 3289 12000
rect 3353 11936 3369 12000
rect 3433 11936 3441 12000
rect 3121 10912 3441 11936
rect 3121 10848 3129 10912
rect 3193 10848 3209 10912
rect 3273 10848 3289 10912
rect 3353 10848 3369 10912
rect 3433 10848 3441 10912
rect 3121 9824 3441 10848
rect 3121 9760 3129 9824
rect 3193 9760 3209 9824
rect 3273 9760 3289 9824
rect 3353 9760 3369 9824
rect 3433 9760 3441 9824
rect 3121 8774 3441 9760
rect 3121 8736 3163 8774
rect 3399 8736 3441 8774
rect 3121 8672 3129 8736
rect 3433 8672 3441 8736
rect 3121 8538 3163 8672
rect 3399 8538 3441 8672
rect 3121 7648 3441 8538
rect 3121 7584 3129 7648
rect 3193 7584 3209 7648
rect 3273 7584 3289 7648
rect 3353 7584 3369 7648
rect 3433 7584 3441 7648
rect 3121 6560 3441 7584
rect 3121 6496 3129 6560
rect 3193 6496 3209 6560
rect 3273 6496 3289 6560
rect 3353 6496 3369 6560
rect 3433 6496 3441 6560
rect 3121 5472 3441 6496
rect 3121 5408 3129 5472
rect 3193 5408 3209 5472
rect 3273 5408 3289 5472
rect 3353 5408 3369 5472
rect 3433 5408 3441 5472
rect 3121 4422 3441 5408
rect 3121 4384 3163 4422
rect 3399 4384 3441 4422
rect 3121 4320 3129 4384
rect 3433 4320 3441 4384
rect 3121 4186 3163 4320
rect 3399 4186 3441 4320
rect 3121 3296 3441 4186
rect 3121 3232 3129 3296
rect 3193 3232 3209 3296
rect 3273 3232 3289 3296
rect 3353 3232 3369 3296
rect 3433 3232 3441 3296
rect 3121 2208 3441 3232
rect 3121 2144 3129 2208
rect 3193 2144 3209 2208
rect 3273 2144 3289 2208
rect 3353 2144 3369 2208
rect 3433 2144 3441 2208
rect 3121 2128 3441 2144
rect 5298 14720 5619 15280
rect 5298 14656 5306 14720
rect 5370 14656 5386 14720
rect 5450 14656 5466 14720
rect 5530 14656 5546 14720
rect 5610 14656 5619 14720
rect 5298 13632 5619 14656
rect 5298 13568 5306 13632
rect 5370 13568 5386 13632
rect 5450 13568 5466 13632
rect 5530 13568 5546 13632
rect 5610 13568 5619 13632
rect 5298 12544 5619 13568
rect 5298 12480 5306 12544
rect 5370 12480 5386 12544
rect 5450 12480 5466 12544
rect 5530 12480 5546 12544
rect 5610 12480 5619 12544
rect 5298 11456 5619 12480
rect 5298 11392 5306 11456
rect 5370 11392 5386 11456
rect 5450 11392 5466 11456
rect 5530 11392 5546 11456
rect 5610 11392 5619 11456
rect 5298 10950 5619 11392
rect 5298 10714 5340 10950
rect 5576 10714 5619 10950
rect 5298 10368 5619 10714
rect 5298 10304 5306 10368
rect 5370 10304 5386 10368
rect 5450 10304 5466 10368
rect 5530 10304 5546 10368
rect 5610 10304 5619 10368
rect 5298 9280 5619 10304
rect 5298 9216 5306 9280
rect 5370 9216 5386 9280
rect 5450 9216 5466 9280
rect 5530 9216 5546 9280
rect 5610 9216 5619 9280
rect 5298 8192 5619 9216
rect 5298 8128 5306 8192
rect 5370 8128 5386 8192
rect 5450 8128 5466 8192
rect 5530 8128 5546 8192
rect 5610 8128 5619 8192
rect 5298 7104 5619 8128
rect 5298 7040 5306 7104
rect 5370 7040 5386 7104
rect 5450 7040 5466 7104
rect 5530 7040 5546 7104
rect 5610 7040 5619 7104
rect 5298 6598 5619 7040
rect 5298 6362 5340 6598
rect 5576 6362 5619 6598
rect 5298 6016 5619 6362
rect 5298 5952 5306 6016
rect 5370 5952 5386 6016
rect 5450 5952 5466 6016
rect 5530 5952 5546 6016
rect 5610 5952 5619 6016
rect 5298 4928 5619 5952
rect 5298 4864 5306 4928
rect 5370 4864 5386 4928
rect 5450 4864 5466 4928
rect 5530 4864 5546 4928
rect 5610 4864 5619 4928
rect 5298 3840 5619 4864
rect 5298 3776 5306 3840
rect 5370 3776 5386 3840
rect 5450 3776 5466 3840
rect 5530 3776 5546 3840
rect 5610 3776 5619 3840
rect 5298 2752 5619 3776
rect 5298 2688 5306 2752
rect 5370 2688 5386 2752
rect 5450 2688 5466 2752
rect 5530 2688 5546 2752
rect 5610 2688 5619 2752
rect 5298 2128 5619 2688
rect 7476 15264 7796 15280
rect 7476 15200 7484 15264
rect 7548 15200 7564 15264
rect 7628 15200 7644 15264
rect 7708 15200 7724 15264
rect 7788 15200 7796 15264
rect 7476 14176 7796 15200
rect 7476 14112 7484 14176
rect 7548 14112 7564 14176
rect 7628 14112 7644 14176
rect 7708 14112 7724 14176
rect 7788 14112 7796 14176
rect 7476 13126 7796 14112
rect 7476 13088 7518 13126
rect 7754 13088 7796 13126
rect 7476 13024 7484 13088
rect 7788 13024 7796 13088
rect 7476 12890 7518 13024
rect 7754 12890 7796 13024
rect 7476 12000 7796 12890
rect 7476 11936 7484 12000
rect 7548 11936 7564 12000
rect 7628 11936 7644 12000
rect 7708 11936 7724 12000
rect 7788 11936 7796 12000
rect 7476 10912 7796 11936
rect 7476 10848 7484 10912
rect 7548 10848 7564 10912
rect 7628 10848 7644 10912
rect 7708 10848 7724 10912
rect 7788 10848 7796 10912
rect 7476 9824 7796 10848
rect 7476 9760 7484 9824
rect 7548 9760 7564 9824
rect 7628 9760 7644 9824
rect 7708 9760 7724 9824
rect 7788 9760 7796 9824
rect 7476 8774 7796 9760
rect 7476 8736 7518 8774
rect 7754 8736 7796 8774
rect 7476 8672 7484 8736
rect 7788 8672 7796 8736
rect 7476 8538 7518 8672
rect 7754 8538 7796 8672
rect 7476 7648 7796 8538
rect 7476 7584 7484 7648
rect 7548 7584 7564 7648
rect 7628 7584 7644 7648
rect 7708 7584 7724 7648
rect 7788 7584 7796 7648
rect 7476 6560 7796 7584
rect 7476 6496 7484 6560
rect 7548 6496 7564 6560
rect 7628 6496 7644 6560
rect 7708 6496 7724 6560
rect 7788 6496 7796 6560
rect 7476 5472 7796 6496
rect 7476 5408 7484 5472
rect 7548 5408 7564 5472
rect 7628 5408 7644 5472
rect 7708 5408 7724 5472
rect 7788 5408 7796 5472
rect 7476 4422 7796 5408
rect 7476 4384 7518 4422
rect 7754 4384 7796 4422
rect 7476 4320 7484 4384
rect 7788 4320 7796 4384
rect 7476 4186 7518 4320
rect 7754 4186 7796 4320
rect 7476 3296 7796 4186
rect 7476 3232 7484 3296
rect 7548 3232 7564 3296
rect 7628 3232 7644 3296
rect 7708 3232 7724 3296
rect 7788 3232 7796 3296
rect 7476 2208 7796 3232
rect 7476 2144 7484 2208
rect 7548 2144 7564 2208
rect 7628 2144 7644 2208
rect 7708 2144 7724 2208
rect 7788 2144 7796 2208
rect 7476 2128 7796 2144
rect 9653 14720 9973 15280
rect 9653 14656 9661 14720
rect 9725 14656 9741 14720
rect 9805 14656 9821 14720
rect 9885 14656 9901 14720
rect 9965 14656 9973 14720
rect 9653 13632 9973 14656
rect 9653 13568 9661 13632
rect 9725 13568 9741 13632
rect 9805 13568 9821 13632
rect 9885 13568 9901 13632
rect 9965 13568 9973 13632
rect 9653 12544 9973 13568
rect 9653 12480 9661 12544
rect 9725 12480 9741 12544
rect 9805 12480 9821 12544
rect 9885 12480 9901 12544
rect 9965 12480 9973 12544
rect 9653 11456 9973 12480
rect 9653 11392 9661 11456
rect 9725 11392 9741 11456
rect 9805 11392 9821 11456
rect 9885 11392 9901 11456
rect 9965 11392 9973 11456
rect 9653 10950 9973 11392
rect 9653 10714 9695 10950
rect 9931 10714 9973 10950
rect 9653 10368 9973 10714
rect 9653 10304 9661 10368
rect 9725 10304 9741 10368
rect 9805 10304 9821 10368
rect 9885 10304 9901 10368
rect 9965 10304 9973 10368
rect 9653 9280 9973 10304
rect 9653 9216 9661 9280
rect 9725 9216 9741 9280
rect 9805 9216 9821 9280
rect 9885 9216 9901 9280
rect 9965 9216 9973 9280
rect 9653 8192 9973 9216
rect 9653 8128 9661 8192
rect 9725 8128 9741 8192
rect 9805 8128 9821 8192
rect 9885 8128 9901 8192
rect 9965 8128 9973 8192
rect 9653 7104 9973 8128
rect 9653 7040 9661 7104
rect 9725 7040 9741 7104
rect 9805 7040 9821 7104
rect 9885 7040 9901 7104
rect 9965 7040 9973 7104
rect 9653 6598 9973 7040
rect 9653 6362 9695 6598
rect 9931 6362 9973 6598
rect 9653 6016 9973 6362
rect 9653 5952 9661 6016
rect 9725 5952 9741 6016
rect 9805 5952 9821 6016
rect 9885 5952 9901 6016
rect 9965 5952 9973 6016
rect 9653 4928 9973 5952
rect 9653 4864 9661 4928
rect 9725 4864 9741 4928
rect 9805 4864 9821 4928
rect 9885 4864 9901 4928
rect 9965 4864 9973 4928
rect 9653 3840 9973 4864
rect 9653 3776 9661 3840
rect 9725 3776 9741 3840
rect 9805 3776 9821 3840
rect 9885 3776 9901 3840
rect 9965 3776 9973 3840
rect 9653 2752 9973 3776
rect 9653 2688 9661 2752
rect 9725 2688 9741 2752
rect 9805 2688 9821 2752
rect 9885 2688 9901 2752
rect 9965 2688 9973 2752
rect 9653 2128 9973 2688
rect 11830 15264 12151 15280
rect 11830 15200 11838 15264
rect 11902 15200 11918 15264
rect 11982 15200 11998 15264
rect 12062 15200 12078 15264
rect 12142 15200 12151 15264
rect 11830 14176 12151 15200
rect 11830 14112 11838 14176
rect 11902 14112 11918 14176
rect 11982 14112 11998 14176
rect 12062 14112 12078 14176
rect 12142 14112 12151 14176
rect 11830 13126 12151 14112
rect 11830 13088 11872 13126
rect 12108 13088 12151 13126
rect 11830 13024 11838 13088
rect 12142 13024 12151 13088
rect 11830 12890 11872 13024
rect 12108 12890 12151 13024
rect 11830 12000 12151 12890
rect 11830 11936 11838 12000
rect 11902 11936 11918 12000
rect 11982 11936 11998 12000
rect 12062 11936 12078 12000
rect 12142 11936 12151 12000
rect 11830 10912 12151 11936
rect 11830 10848 11838 10912
rect 11902 10848 11918 10912
rect 11982 10848 11998 10912
rect 12062 10848 12078 10912
rect 12142 10848 12151 10912
rect 11830 9824 12151 10848
rect 11830 9760 11838 9824
rect 11902 9760 11918 9824
rect 11982 9760 11998 9824
rect 12062 9760 12078 9824
rect 12142 9760 12151 9824
rect 11830 8774 12151 9760
rect 11830 8736 11872 8774
rect 12108 8736 12151 8774
rect 11830 8672 11838 8736
rect 12142 8672 12151 8736
rect 11830 8538 11872 8672
rect 12108 8538 12151 8672
rect 11830 7648 12151 8538
rect 11830 7584 11838 7648
rect 11902 7584 11918 7648
rect 11982 7584 11998 7648
rect 12062 7584 12078 7648
rect 12142 7584 12151 7648
rect 11830 6560 12151 7584
rect 11830 6496 11838 6560
rect 11902 6496 11918 6560
rect 11982 6496 11998 6560
rect 12062 6496 12078 6560
rect 12142 6496 12151 6560
rect 11830 5472 12151 6496
rect 11830 5408 11838 5472
rect 11902 5408 11918 5472
rect 11982 5408 11998 5472
rect 12062 5408 12078 5472
rect 12142 5408 12151 5472
rect 11830 4422 12151 5408
rect 11830 4384 11872 4422
rect 12108 4384 12151 4422
rect 11830 4320 11838 4384
rect 12142 4320 12151 4384
rect 11830 4186 11872 4320
rect 12108 4186 12151 4320
rect 11830 3296 12151 4186
rect 11830 3232 11838 3296
rect 11902 3232 11918 3296
rect 11982 3232 11998 3296
rect 12062 3232 12078 3296
rect 12142 3232 12151 3296
rect 11830 2208 12151 3232
rect 11830 2144 11838 2208
rect 11902 2144 11918 2208
rect 11982 2144 11998 2208
rect 12062 2144 12078 2208
rect 12142 2144 12151 2208
rect 11830 2128 12151 2144
<< via4 >>
rect 3163 13088 3399 13126
rect 3163 13024 3193 13088
rect 3193 13024 3209 13088
rect 3209 13024 3273 13088
rect 3273 13024 3289 13088
rect 3289 13024 3353 13088
rect 3353 13024 3369 13088
rect 3369 13024 3399 13088
rect 3163 12890 3399 13024
rect 3163 8736 3399 8774
rect 3163 8672 3193 8736
rect 3193 8672 3209 8736
rect 3209 8672 3273 8736
rect 3273 8672 3289 8736
rect 3289 8672 3353 8736
rect 3353 8672 3369 8736
rect 3369 8672 3399 8736
rect 3163 8538 3399 8672
rect 3163 4384 3399 4422
rect 3163 4320 3193 4384
rect 3193 4320 3209 4384
rect 3209 4320 3273 4384
rect 3273 4320 3289 4384
rect 3289 4320 3353 4384
rect 3353 4320 3369 4384
rect 3369 4320 3399 4384
rect 3163 4186 3399 4320
rect 5340 10714 5576 10950
rect 5340 6362 5576 6598
rect 7518 13088 7754 13126
rect 7518 13024 7548 13088
rect 7548 13024 7564 13088
rect 7564 13024 7628 13088
rect 7628 13024 7644 13088
rect 7644 13024 7708 13088
rect 7708 13024 7724 13088
rect 7724 13024 7754 13088
rect 7518 12890 7754 13024
rect 7518 8736 7754 8774
rect 7518 8672 7548 8736
rect 7548 8672 7564 8736
rect 7564 8672 7628 8736
rect 7628 8672 7644 8736
rect 7644 8672 7708 8736
rect 7708 8672 7724 8736
rect 7724 8672 7754 8736
rect 7518 8538 7754 8672
rect 7518 4384 7754 4422
rect 7518 4320 7548 4384
rect 7548 4320 7564 4384
rect 7564 4320 7628 4384
rect 7628 4320 7644 4384
rect 7644 4320 7708 4384
rect 7708 4320 7724 4384
rect 7724 4320 7754 4384
rect 7518 4186 7754 4320
rect 9695 10714 9931 10950
rect 9695 6362 9931 6598
rect 11872 13088 12108 13126
rect 11872 13024 11902 13088
rect 11902 13024 11918 13088
rect 11918 13024 11982 13088
rect 11982 13024 11998 13088
rect 11998 13024 12062 13088
rect 12062 13024 12078 13088
rect 12078 13024 12108 13088
rect 11872 12890 12108 13024
rect 11872 8736 12108 8774
rect 11872 8672 11902 8736
rect 11902 8672 11918 8736
rect 11918 8672 11982 8736
rect 11982 8672 11998 8736
rect 11998 8672 12062 8736
rect 12062 8672 12078 8736
rect 12078 8672 12108 8736
rect 11872 8538 12108 8672
rect 11872 4384 12108 4422
rect 11872 4320 11902 4384
rect 11902 4320 11918 4384
rect 11918 4320 11982 4384
rect 11982 4320 11998 4384
rect 11998 4320 12062 4384
rect 12062 4320 12078 4384
rect 12078 4320 12108 4384
rect 11872 4186 12108 4320
<< metal5 >>
rect 1104 13126 14168 13168
rect 1104 12890 3163 13126
rect 3399 12890 7518 13126
rect 7754 12890 11872 13126
rect 12108 12890 14168 13126
rect 1104 12848 14168 12890
rect 1104 10950 14168 10992
rect 1104 10714 5340 10950
rect 5576 10714 9695 10950
rect 9931 10714 14168 10950
rect 1104 10672 14168 10714
rect 1104 8774 14168 8816
rect 1104 8538 3163 8774
rect 3399 8538 7518 8774
rect 7754 8538 11872 8774
rect 12108 8538 14168 8774
rect 1104 8496 14168 8538
rect 1104 6598 14168 6640
rect 1104 6362 5340 6598
rect 5576 6362 9695 6598
rect 9931 6362 14168 6598
rect 1104 6320 14168 6362
rect 1104 4422 14168 4464
rect 1104 4186 3163 4422
rect 3399 4186 7518 4422
rect 7754 4186 11872 4422
rect 12108 4186 14168 4422
rect 1104 4144 14168 4186
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1619150647
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform -1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 2116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1619150647
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1619150647
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 3220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1619150647
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1619150647
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1619150647
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1619150647
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1619150647
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1619150647
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1619150647
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1619150647
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51
timestamp 1619150647
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1619150647
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform -1 0 9384 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1619150647
transform -1 0 8188 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 8188 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1619150647
transform 1 0 7544 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _25_
timestamp 1619150647
transform 1 0 9752 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1619150647
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1619150647
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1619150647
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1619150647
transform 1 0 10304 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1619150647
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1619150647
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1619150647
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1619150647
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1619150647
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1619150647
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1619150647
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1619150647
transform -1 0 14168 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1619150647
transform -1 0 14168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output2
timestamp 1619150647
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1619150647
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1619150647
transform 1 0 13524 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1619150647
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1619150647
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1619150647
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1619150647
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1619150647
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1619150647
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1619150647
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1619150647
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1619150647
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 8096 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_66
timestamp 1619150647
transform 1 0 7176 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1619150647
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_79
timestamp 1619150647
transform 1 0 8372 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 10672 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 9752 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1619150647
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_87
timestamp 1619150647
transform 1 0 9108 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1619150647
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_100
timestamp 1619150647
transform 1 0 10304 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_107
timestamp 1619150647
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_119
timestamp 1619150647
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1619150647
transform -1 0 14168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_131
timestamp 1619150647
transform 1 0 13156 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1619150647
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1619150647
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1619150647
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1619150647
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1619150647
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1619150647
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1619150647
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1619150647
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1619150647
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1619150647
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1619150647
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1619150647
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1619150647
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1619150647
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1619150647
transform -1 0 14168 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1619150647
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1619150647
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1619150647
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1619150647
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1619150647
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1619150647
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1619150647
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1619150647
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1619150647
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1619150647
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1619150647
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1619150647
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform -1 0 9752 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1619150647
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_94
timestamp 1619150647
transform 1 0 9752 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_106
timestamp 1619150647
transform 1 0 10856 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_118
timestamp 1619150647
transform 1 0 11960 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1619150647
transform -1 0 14168 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_130
timestamp 1619150647
transform 1 0 13064 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_138
timestamp 1619150647
transform 1 0 13800 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1619150647
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1619150647
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1619150647
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1619150647
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1619150647
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1619150647
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1619150647
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1619150647
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1619150647
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1619150647
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1619150647
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1619150647
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1619150647
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1619150647
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1619150647
transform -1 0 14168 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1619150647
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1619150647
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1619150647
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1619150647
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1619150647
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1619150647
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1619150647
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1619150647
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1619150647
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1619150647
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1619150647
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1619150647
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1619150647
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1619150647
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1619150647
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1619150647
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1619150647
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1619150647
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1619150647
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1619150647
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1619150647
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1619150647
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1619150647
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1619150647
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1619150647
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1619150647
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1619150647
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1619150647
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1619150647
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1619150647
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1619150647
transform -1 0 14168 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1619150647
transform -1 0 14168 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1619150647
transform 1 0 13524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1619150647
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1619150647
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1619150647
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1619150647
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1619150647
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1619150647
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1619150647
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1619150647
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1619150647
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1619150647
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1619150647
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1619150647
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1619150647
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1619150647
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1619150647
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1619150647
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1619150647
transform -1 0 14168 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1619150647
transform 1 0 13524 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1619150647
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1619150647
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1619150647
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1619150647
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1619150647
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1619150647
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1619150647
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1619150647
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform -1 0 10304 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_9_70
timestamp 1619150647
transform 1 0 7544 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1619150647
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_100
timestamp 1619150647
transform 1 0 10304 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1619150647
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1619150647
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1619150647
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1619150647
transform -1 0 14168 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1619150647
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1619150647
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1619150647
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1619150647
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1619150647
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1619150647
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1619150647
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1619150647
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1619150647
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1619150647
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1619150647
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1619150647
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1619150647
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1619150647
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1619150647
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1619150647
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1619150647
transform -1 0 14168 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1619150647
transform 1 0 13524 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1619150647
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1619150647
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1619150647
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1619150647
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1619150647
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1619150647
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1619150647
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1619150647
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1619150647
transform 1 0 8556 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_70
timestamp 1619150647
transform 1 0 7544 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_78
timestamp 1619150647
transform 1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_84
timestamp 1619150647
transform 1 0 8832 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_96
timestamp 1619150647
transform 1 0 9936 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1619150647
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_108
timestamp 1619150647
transform 1 0 11040 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1619150647
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1619150647
transform -1 0 14168 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1619150647
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1619150647
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1619150647
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1619150647
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1619150647
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1619150647
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1619150647
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1619150647
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1619150647
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _21_
timestamp 1619150647
transform -1 0 8188 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_66
timestamp 1619150647
transform 1 0 7176 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_77
timestamp 1619150647
transform 1 0 8188 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _14_
timestamp 1619150647
transform -1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1619150647
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1619150647
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_87
timestamp 1619150647
transform 1 0 9108 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_95
timestamp 1619150647
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_100
timestamp 1619150647
transform 1 0 10304 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_112
timestamp 1619150647
transform 1 0 11408 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_124
timestamp 1619150647
transform 1 0 12512 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1619150647
transform -1 0 14168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_136
timestamp 1619150647
transform 1 0 13616 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1619150647
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1619150647
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1619150647
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1619150647
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1619150647
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1619150647
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1619150647
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1619150647
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1619150647
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1619150647
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1619150647
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _20_
timestamp 1619150647
transform -1 0 6716 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _29_
timestamp 1619150647
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1619150647
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1619150647
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_58
timestamp 1619150647
transform 1 0 6440 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1619150647
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_54
timestamp 1619150647
transform 1 0 6072 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1619150647
transform 1 0 6716 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _19_
timestamp 1619150647
transform -1 0 8464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 7084 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_78
timestamp 1619150647
transform 1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_73
timestamp 1619150647
transform 1 0 7820 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_80
timestamp 1619150647
transform 1 0 8464 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_87
timestamp 1619150647
transform 1 0 9108 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1619150647
transform 1 0 9476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1619150647
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1619150647
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform -1 0 9476 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_95
timestamp 1619150647
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1619150647
transform 1 0 10672 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_95
timestamp 1619150647
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform -1 0 10672 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _26_
timestamp 1619150647
transform 1 0 10028 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1619150647
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1619150647
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1619150647
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_113
timestamp 1619150647
transform 1 0 11500 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_125
timestamp 1619150647
transform 1 0 12604 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1619150647
transform -1 0 14168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1619150647
transform -1 0 14168 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1619150647
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_137
timestamp 1619150647
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1619150647
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1619150647
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1619150647
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1619150647
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1619150647
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _28_
timestamp 1619150647
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1619150647
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1619150647
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_58
timestamp 1619150647
transform 1 0 6440 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_78
timestamp 1619150647
transform 1 0 8280 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _27_
timestamp 1619150647
transform 1 0 8924 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_84
timestamp 1619150647
transform 1 0 8832 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1619150647
transform 1 0 10396 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform 1 0 10764 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1619150647
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_109
timestamp 1619150647
transform 1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1619150647
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1619150647
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1619150647
transform -1 0 14168 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1619150647
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1619150647
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output4
timestamp 1619150647
transform -1 0 2116 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1619150647
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_11
timestamp 1619150647
transform 1 0 2116 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1619150647
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_23
timestamp 1619150647
transform 1 0 3220 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1619150647
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1619150647
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1619150647
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1619150647
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1619150647
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _16_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1619150647
transform -1 0 9936 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1619150647
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1619150647
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_96
timestamp 1619150647
transform 1 0 9936 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_108
timestamp 1619150647
transform 1 0 11040 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_120
timestamp 1619150647
transform 1 0 12144 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1619150647
transform -1 0 14168 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_132
timestamp 1619150647
transform 1 0 13248 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_138
timestamp 1619150647
transform 1 0 13800 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1619150647
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1619150647
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1619150647
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1619150647
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1619150647
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1619150647
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1619150647
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1619150647
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1619150647
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1619150647
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1619150647
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1619150647
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1619150647
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1619150647
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1619150647
transform -1 0 14168 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output3
timestamp 1619150647
transform 1 0 13156 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1619150647
transform 1 0 12788 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1619150647
transform 1 0 13524 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1619150647
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1619150647
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1619150647
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1619150647
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1619150647
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1619150647
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1619150647
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1619150647
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1619150647
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1619150647
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1619150647
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1619150647
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1619150647
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1619150647
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1619150647
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1619150647
transform -1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1619150647
transform 1 0 13524 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1619150647
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1619150647
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1619150647
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1619150647
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1619150647
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1619150647
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1619150647
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1619150647
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1619150647
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1619150647
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1619150647
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1619150647
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1619150647
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1619150647
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1619150647
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1619150647
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1619150647
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1619150647
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1619150647
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1619150647
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1619150647
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1619150647
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1619150647
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1619150647
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1619150647
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1619150647
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1619150647
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1619150647
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1619150647
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1619150647
transform -1 0 14168 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1619150647
transform -1 0 14168 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1619150647
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1619150647
transform 1 0 13524 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1619150647
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1619150647
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1619150647
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1619150647
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1619150647
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1619150647
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1619150647
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1619150647
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1619150647
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1619150647
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1619150647
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1619150647
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1619150647
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1619150647
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1619150647
transform -1 0 14168 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1619150647
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1619150647
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1619150647
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1619150647
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1619150647
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1619150647
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1619150647
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1619150647
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1619150647
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1619150647
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1619150647
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1619150647
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1619150647
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1619150647
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1619150647
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1619150647
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1619150647
transform -1 0 14168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1619150647
transform 1 0 13524 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1619150647
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1619150647
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1619150647
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1619150647
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1619150647
transform -1 0 4600 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1619150647
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1619150647
transform 1 0 3864 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_38
timestamp 1619150647
transform 1 0 4600 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1619150647
transform 1 0 6440 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_50
timestamp 1619150647
transform 1 0 5704 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_59
timestamp 1619150647
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_71
timestamp 1619150647
transform 1 0 7636 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1619150647
transform 1 0 8740 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1619150647
transform 1 0 9108 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_88
timestamp 1619150647
transform 1 0 9200 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_100
timestamp 1619150647
transform 1 0 10304 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1619150647
transform 1 0 11776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_112
timestamp 1619150647
transform 1 0 11408 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_117
timestamp 1619150647
transform 1 0 11868 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1619150647
transform -1 0 14168 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_129
timestamp 1619150647
transform 1 0 12972 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1619150647
transform 1 0 13708 0 1 14688
box -38 -48 222 592
<< labels >>
rlabel metal2 s 11058 16635 11114 17435 6 clk
port 0 nsew signal input
rlabel metal2 s 478 0 534 800 6 counter[0]
port 1 nsew signal tristate
rlabel metal3 s 14491 688 15291 808 6 counter[1]
port 2 nsew signal tristate
rlabel metal3 s 14491 11568 15291 11688 6 counter[2]
port 3 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 counter[3]
port 4 nsew signal tristate
rlabel metal2 s 3698 16635 3754 17435 6 counter[4]
port 5 nsew signal tristate
rlabel metal2 s 7838 0 7894 800 6 counter[5]
port 6 nsew signal tristate
rlabel metal4 s 11831 2128 12151 15280 6 VPWR
port 7 nsew power bidirectional
rlabel metal4 s 7476 2128 7796 15280 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 3121 2128 3441 15280 6 VPWR
port 9 nsew power bidirectional
rlabel metal5 s 1104 12848 14168 13168 6 VPWR
port 10 nsew power bidirectional
rlabel metal5 s 1104 8496 14168 8816 6 VPWR
port 11 nsew power bidirectional
rlabel metal5 s 1104 4144 14168 4464 6 VPWR
port 12 nsew power bidirectional
rlabel metal4 s 9653 2128 9973 15280 6 VGND
port 13 nsew ground bidirectional
rlabel metal4 s 5299 2128 5619 15280 6 VGND
port 14 nsew ground bidirectional
rlabel metal5 s 1104 10672 14168 10992 6 VGND
port 15 nsew ground bidirectional
rlabel metal5 s 1104 6320 14168 6640 6 VGND
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15291 17435
<< end >>
