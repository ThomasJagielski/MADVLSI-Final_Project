magic
tech sky130A
timestamp 1620755988
<< nwell >>
rect -135 35 1195 375
<< pmos >>
rect 5 55 65 355
rect 215 55 275 355
rect 335 55 395 355
rect 455 55 515 355
rect 575 55 635 355
rect 695 55 755 355
rect 815 55 875 355
rect 935 55 995 355
rect 1055 55 1115 355
<< pdiff >>
rect -55 340 5 355
rect -55 70 -40 340
rect -10 70 5 340
rect -55 55 5 70
rect 65 340 125 355
rect 65 70 80 340
rect 110 70 125 340
rect 65 55 125 70
rect 155 340 215 355
rect 155 70 170 340
rect 200 70 215 340
rect 155 55 215 70
rect 275 340 335 355
rect 275 70 290 340
rect 320 70 335 340
rect 275 55 335 70
rect 395 340 455 355
rect 395 70 410 340
rect 440 70 455 340
rect 395 55 455 70
rect 515 340 575 355
rect 515 70 530 340
rect 560 70 575 340
rect 515 55 575 70
rect 635 340 695 355
rect 635 70 650 340
rect 680 70 695 340
rect 635 55 695 70
rect 755 340 815 355
rect 755 70 770 340
rect 800 70 815 340
rect 755 55 815 70
rect 875 340 935 355
rect 875 70 890 340
rect 920 70 935 340
rect 875 55 935 70
rect 995 340 1055 355
rect 995 70 1010 340
rect 1040 70 1055 340
rect 995 55 1055 70
rect 1115 340 1175 355
rect 1115 70 1130 340
rect 1160 70 1175 340
rect 1115 55 1175 70
<< pdiffc >>
rect -40 70 -10 340
rect 80 70 110 340
rect 170 70 200 340
rect 290 70 320 340
rect 410 70 440 340
rect 530 70 560 340
rect 650 70 680 340
rect 770 70 800 340
rect 890 70 920 340
rect 1010 70 1040 340
rect 1130 70 1160 340
<< nsubdiff >>
rect -115 340 -55 355
rect -115 70 -100 340
rect -70 70 -55 340
rect -115 55 -55 70
<< nsubdiffcont >>
rect -100 70 -70 340
<< poly >>
rect 5 355 65 370
rect 215 355 275 370
rect 335 355 395 370
rect 455 355 515 370
rect 575 355 635 370
rect 695 355 755 370
rect 815 355 875 370
rect 935 355 995 370
rect 1055 355 1115 370
rect 5 45 65 55
rect 215 45 275 55
rect 335 45 395 55
rect 455 45 515 55
rect 575 45 635 55
rect 695 45 755 55
rect 815 45 875 55
rect 935 45 995 55
rect 1055 45 1115 55
rect 5 30 1115 45
<< locali >>
rect 280 370 1050 390
rect -110 340 0 350
rect -110 70 -100 340
rect -70 70 -40 340
rect -10 70 0 340
rect -110 60 0 70
rect 70 340 120 350
rect 70 70 80 340
rect 110 70 120 340
rect 70 60 120 70
rect 160 340 210 350
rect 160 70 170 340
rect 200 70 210 340
rect 160 60 210 70
rect 280 340 330 370
rect 280 70 290 340
rect 320 70 330 340
rect 280 60 330 70
rect 400 340 450 350
rect 400 70 410 340
rect 440 70 450 340
rect 400 60 450 70
rect 520 340 570 370
rect 520 70 530 340
rect 560 70 570 340
rect 520 60 570 70
rect 640 340 690 350
rect 640 70 650 340
rect 680 70 690 340
rect 640 60 690 70
rect 760 340 810 370
rect 760 70 770 340
rect 800 70 810 340
rect 760 60 810 70
rect 880 340 930 350
rect 880 70 890 340
rect 920 70 930 340
rect 880 60 930 70
rect 1000 340 1050 370
rect 1000 70 1010 340
rect 1040 70 1050 340
rect 1000 60 1050 70
rect 1120 340 1170 350
rect 1120 70 1130 340
rect 1160 70 1170 340
rect 1120 60 1170 70
<< viali >>
rect -100 70 -70 340
rect -40 70 -10 340
rect 170 70 200 340
rect 410 70 440 340
rect 650 70 680 340
rect 890 70 920 340
rect 1130 70 1160 340
<< metal1 >>
rect -115 340 1175 350
rect -115 70 -100 340
rect -70 70 -40 340
rect -10 70 170 340
rect 200 70 410 340
rect 440 70 650 340
rect 680 70 890 340
rect 920 70 1130 340
rect 1160 70 1175 340
rect -115 60 1175 70
<< end >>
