magic
tech sky130A
timestamp 1620747333
<< poly >>
rect 8780 1505 8825 1515
rect 8780 1485 8790 1505
rect 8815 1485 8825 1505
rect 8780 1475 8825 1485
rect 8780 -1760 8825 -1750
rect 8780 -1780 8790 -1760
rect 8815 -1780 8825 -1760
rect 8780 -1790 8825 -1780
rect -85 -2000 -35 -1985
rect -85 -2020 -70 -2000
rect -50 -2020 -35 -2000
rect -85 -2125 -35 -2020
rect -85 -2145 -70 -2125
rect -50 -2145 -35 -2125
rect -85 -2160 -35 -2145
<< polycont >>
rect 8790 1485 8815 1505
rect 8790 -1780 8815 -1760
rect -70 -2020 -50 -2000
rect -70 -2145 -50 -2125
<< locali >>
rect -165 3390 55 3425
rect -165 -2055 -135 3390
rect -75 3000 35 3040
rect -75 -1985 -45 3000
rect 8780 1505 8825 1515
rect 8780 1485 8790 1505
rect 8815 1485 8825 1505
rect 8780 1475 8825 1485
rect 8980 1285 9085 1305
rect 8980 1215 9000 1285
rect 9065 1215 9085 1285
rect 8980 1180 9085 1215
rect 7345 1140 9085 1180
rect 8980 -385 9085 1140
rect 8980 -405 9260 -385
rect 8780 -1760 8825 -1750
rect 8780 -1780 8790 -1760
rect 8815 -1780 8825 -1760
rect 8780 -1790 8825 -1780
rect -85 -2000 -35 -1985
rect -85 -2020 -70 -2000
rect -50 -2020 -35 -2000
rect -85 -2035 -35 -2020
rect -165 -2090 65 -2055
rect -85 -2125 -35 -2110
rect -85 -2145 -70 -2125
rect -50 -2145 -35 -2125
rect -85 -2440 -35 -2145
rect -85 -2480 50 -2440
rect 8980 -3920 9085 -3900
rect 8980 -3990 9000 -3920
rect 9065 -3990 9085 -3920
rect 8980 -4300 9085 -3990
rect 7365 -4340 9085 -4300
<< viali >>
rect 8790 1485 8815 1505
rect 9000 1215 9065 1285
rect 8790 -1780 8815 -1760
rect 9000 -3990 9065 -3920
<< metal1 >>
rect -235 3285 35 3325
rect -235 -2785 -200 3285
rect 8780 1510 8825 1515
rect 8780 1480 8785 1510
rect 8820 1480 8825 1510
rect 8780 1455 8825 1480
rect 7440 1435 8825 1455
rect 7440 1090 7460 1435
rect 7240 1070 7460 1090
rect 6220 205 6770 930
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 6220 110 6770 120
rect -120 -5 25 15
rect -120 -2155 -75 -5
rect 6220 -90 6770 -80
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -970 6770 -175
rect 5335 -1505 6770 -970
rect 8780 -100 8825 1435
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 8780 -135 10025 -100
rect 5335 -1975 5645 -1505
rect 8780 -1755 8825 -135
rect 8780 -1785 8785 -1755
rect 8820 -1785 8825 -1755
rect 8780 -1790 8825 -1785
rect 8780 -1885 8825 -1825
rect -120 -2195 45 -2155
rect 4625 -2285 5645 -1975
rect 4625 -2405 4725 -2285
rect 5545 -2405 5645 -2285
rect -235 -2820 25 -2785
rect 8990 -3920 9075 -3910
rect 8990 -3990 9000 -3920
rect 9065 -3990 9075 -3920
rect 8990 -4000 9075 -3990
<< via1 >>
rect 8785 1505 8820 1510
rect 8785 1485 8790 1505
rect 8790 1485 8815 1505
rect 8815 1485 8820 1505
rect 8785 1480 8820 1485
rect 6230 120 6760 205
rect 6230 -175 6760 -90
rect 9000 1215 9065 1285
rect 8785 -1760 8820 -1755
rect 8785 -1780 8790 -1760
rect 8790 -1780 8815 -1760
rect 8815 -1780 8820 -1760
rect 8785 -1785 8820 -1780
rect 9000 -3990 9065 -3920
<< metal2 >>
rect -235 2720 15 2760
rect -235 -3350 -200 2720
rect 8780 1510 8825 1515
rect 8780 1480 8785 1510
rect 8820 1480 8825 1510
rect 8780 1475 8825 1480
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 4005 685 4425 835
rect 4005 470 4270 685
rect 4005 405 4015 470
rect 4260 405 4270 470
rect 4005 395 4270 405
rect 6220 205 6770 215
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 6220 110 6770 120
rect -120 -5 25 15
rect -120 -2720 -75 -5
rect 4025 -65 4355 -55
rect 4025 -145 4035 -65
rect 4345 -145 4355 -65
rect 4025 -2405 4355 -145
rect 6220 -90 6770 -80
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -185 6770 -175
rect 8780 -1755 8825 -1750
rect 8780 -1785 8785 -1755
rect 8820 -1785 8825 -1755
rect 8780 -1790 8825 -1785
rect -120 -2760 30 -2720
rect -235 -3390 60 -3350
rect 8990 -3920 9075 -3910
rect 8990 -3990 9000 -3920
rect 9065 -3990 9075 -3920
rect 8990 -4000 9075 -3990
<< via2 >>
rect 8785 1480 8820 1510
rect 9000 1215 9065 1285
rect 4015 405 4260 470
rect 6230 120 6760 205
rect 4035 -145 4345 -65
rect 6230 -175 6760 -90
rect 8785 -1785 8820 -1755
rect 9000 -3990 9065 -3920
<< metal3 >>
rect -250 3155 1405 3210
rect -250 -2270 -190 3155
rect 8775 1510 8830 1585
rect 8775 1480 8785 1510
rect 8820 1480 8830 1510
rect 8775 1475 8830 1480
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 4005 470 4270 480
rect 4005 405 4015 470
rect 4260 405 4270 470
rect 4005 395 4270 405
rect 4025 -55 4270 395
rect 6220 205 6770 215
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 4025 -65 4355 -55
rect 4025 -145 4035 -65
rect 4345 -145 4355 -65
rect 4025 -155 4355 -145
rect 6220 -90 6770 120
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -185 6770 -175
rect 8775 -1755 8830 -1750
rect 8775 -1785 8785 -1755
rect 8820 -1785 8830 -1755
rect 8775 -1855 8830 -1785
rect -255 -2320 1260 -2270
rect 8990 -3920 9075 -3910
rect 8990 -3990 9000 -3920
rect 9065 -3990 9075 -3920
rect 8990 -4000 9075 -3990
<< via3 >>
rect 9000 1215 9065 1285
rect 9000 -3990 9065 -3920
<< metal4 >>
rect 8980 1285 9085 1840
rect 8980 1215 9000 1285
rect 9065 1215 9085 1285
rect 8980 -2125 9085 1215
rect 8980 -3920 9085 -3320
rect 8980 -3990 9000 -3920
rect 9065 -3990 9085 -3920
rect 8980 -4065 9085 -3990
use middle_ping_pong_amplifier  middle_ping_pong_amplifier_0
timestamp 1620710927
transform 1 0 12905 0 1 -1890
box -3700 -30 4680 3175
use cap8to1  cap8to1_0
timestamp 1620746045
transform 1 0 8760 0 1 -3670
box 5 30 3785 1860
use cap8to1  cap8to1_1
timestamp 1620746045
transform 1 0 8760 0 1 1495
box 5 30 3785 1860
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_0
timestamp 1620746045
transform 1 0 3930 0 1 570
box -3935 -575 4700 4735
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_1
timestamp 1620746045
transform 1 0 3950 0 1 -4910
box -3935 -575 4700 4735
<< end >>
