magic
tech sky130A
timestamp 1620532465
<< nwell >>
rect -205 4600 2065 4800
rect 330 4480 435 4600
rect 1510 4490 1615 4600
rect -205 3875 2065 4075
rect 340 3765 445 3875
rect 1420 3755 1525 3875
rect -205 2940 2065 3140
rect 215 2745 375 2940
rect 1605 2745 1765 2940
<< nmos >>
rect -120 4295 -60 4445
rect 0 4295 60 4445
rect 120 4295 180 4445
rect 240 4295 300 4445
rect 360 4295 420 4445
rect 480 4295 540 4445
rect 600 4295 660 4445
rect 720 4295 780 4445
rect 840 4295 900 4445
rect 960 4295 1020 4445
rect 1080 4295 1140 4445
rect 1200 4295 1260 4445
rect 1320 4295 1380 4445
rect 1440 4295 1500 4445
rect 1560 4295 1620 4445
rect 1680 4295 1740 4445
rect 1800 4295 1860 4445
rect 1920 4295 1980 4445
rect -120 3460 -60 3610
rect 0 3460 60 3610
rect 120 3460 180 3610
rect 240 3460 300 3610
rect 360 3460 420 3610
rect 480 3460 540 3610
rect 600 3460 660 3610
rect 720 3460 780 3610
rect 840 3460 900 3610
rect 960 3460 1020 3610
rect 1080 3460 1140 3610
rect 1200 3460 1260 3610
rect 1320 3460 1380 3610
rect 1440 3460 1500 3610
rect 1560 3460 1620 3610
rect 1680 3460 1740 3610
rect 1800 3460 1860 3610
rect 1920 3460 1980 3610
rect -120 2430 -60 2580
rect 0 2430 60 2580
rect 120 2430 180 2580
rect 240 2430 300 2580
rect 360 2430 420 2580
rect 480 2430 540 2580
rect 600 2430 660 2580
rect 720 2430 780 2580
rect 840 2430 900 2580
rect 960 2430 1020 2580
rect 1080 2430 1140 2580
rect 1200 2430 1260 2580
rect 1320 2430 1380 2580
rect 1440 2430 1500 2580
rect 1560 2430 1620 2580
rect 1680 2430 1740 2580
rect 1800 2430 1860 2580
rect 1920 2430 1980 2580
<< pmos >>
rect -120 4625 -60 4775
rect 0 4625 60 4775
rect 120 4625 180 4775
rect 240 4625 300 4775
rect 360 4625 420 4775
rect 480 4625 540 4775
rect 600 4625 660 4775
rect 720 4625 780 4775
rect 840 4625 900 4775
rect 960 4625 1020 4775
rect 1080 4625 1140 4775
rect 1200 4625 1260 4775
rect 1320 4625 1380 4775
rect 1440 4625 1500 4775
rect 1560 4625 1620 4775
rect 1680 4625 1740 4775
rect 1800 4625 1860 4775
rect 1920 4625 1980 4775
rect -120 3900 -60 4050
rect 0 3900 60 4050
rect 120 3900 180 4050
rect 240 3900 300 4050
rect 360 3900 420 4050
rect 480 3900 540 4050
rect 600 3900 660 4050
rect 720 3900 780 4050
rect 840 3900 900 4050
rect 960 3900 1020 4050
rect 1080 3900 1140 4050
rect 1200 3900 1260 4050
rect 1320 3900 1380 4050
rect 1440 3900 1500 4050
rect 1560 3900 1620 4050
rect 1680 3900 1740 4050
rect 1800 3900 1860 4050
rect 1920 3900 1980 4050
rect -120 2965 -60 3115
rect 0 2965 60 3115
rect 120 2965 180 3115
rect 240 2965 300 3115
rect 360 2965 420 3115
rect 480 2965 540 3115
rect 600 2965 660 3115
rect 720 2965 780 3115
rect 840 2965 900 3115
rect 960 2965 1020 3115
rect 1080 2965 1140 3115
rect 1200 2965 1260 3115
rect 1320 2965 1380 3115
rect 1440 2965 1500 3115
rect 1560 2965 1620 3115
rect 1680 2965 1740 3115
rect 1800 2965 1860 3115
rect 1920 2965 1980 3115
<< ndiff >>
rect -180 4430 -120 4445
rect -180 4310 -165 4430
rect -135 4310 -120 4430
rect -180 4295 -120 4310
rect -60 4430 0 4445
rect -60 4310 -45 4430
rect -15 4310 0 4430
rect -60 4295 0 4310
rect 60 4430 120 4445
rect 60 4310 75 4430
rect 105 4310 120 4430
rect 60 4295 120 4310
rect 180 4430 240 4445
rect 180 4310 195 4430
rect 225 4310 240 4430
rect 180 4295 240 4310
rect 300 4430 360 4445
rect 300 4310 315 4430
rect 345 4310 360 4430
rect 300 4295 360 4310
rect 420 4430 480 4445
rect 420 4310 435 4430
rect 465 4310 480 4430
rect 420 4295 480 4310
rect 540 4430 600 4445
rect 540 4310 555 4430
rect 585 4310 600 4430
rect 540 4295 600 4310
rect 660 4430 720 4445
rect 660 4310 675 4430
rect 705 4310 720 4430
rect 660 4295 720 4310
rect 780 4430 840 4445
rect 780 4310 795 4430
rect 825 4310 840 4430
rect 780 4295 840 4310
rect 900 4430 960 4445
rect 900 4310 915 4430
rect 945 4310 960 4430
rect 900 4295 960 4310
rect 1020 4430 1080 4445
rect 1020 4310 1035 4430
rect 1065 4310 1080 4430
rect 1020 4295 1080 4310
rect 1140 4430 1200 4445
rect 1140 4310 1155 4430
rect 1185 4310 1200 4430
rect 1140 4295 1200 4310
rect 1260 4430 1320 4445
rect 1260 4310 1275 4430
rect 1305 4310 1320 4430
rect 1260 4295 1320 4310
rect 1380 4430 1440 4445
rect 1380 4310 1395 4430
rect 1425 4310 1440 4430
rect 1380 4295 1440 4310
rect 1500 4430 1560 4445
rect 1500 4310 1515 4430
rect 1545 4310 1560 4430
rect 1500 4295 1560 4310
rect 1620 4430 1680 4445
rect 1620 4310 1635 4430
rect 1665 4310 1680 4430
rect 1620 4295 1680 4310
rect 1740 4430 1800 4445
rect 1740 4310 1755 4430
rect 1785 4310 1800 4430
rect 1740 4295 1800 4310
rect 1860 4430 1920 4445
rect 1860 4310 1875 4430
rect 1905 4310 1920 4430
rect 1860 4295 1920 4310
rect 1980 4430 2040 4445
rect 1980 4310 1995 4430
rect 2025 4310 2040 4430
rect 1980 4295 2040 4310
rect -180 3595 -120 3610
rect -180 3475 -165 3595
rect -135 3475 -120 3595
rect -180 3460 -120 3475
rect -60 3595 0 3610
rect -60 3475 -45 3595
rect -15 3475 0 3595
rect -60 3460 0 3475
rect 60 3595 120 3610
rect 60 3475 75 3595
rect 105 3475 120 3595
rect 60 3460 120 3475
rect 180 3595 240 3610
rect 180 3475 195 3595
rect 225 3475 240 3595
rect 180 3460 240 3475
rect 300 3595 360 3610
rect 300 3475 315 3595
rect 345 3475 360 3595
rect 300 3460 360 3475
rect 420 3595 480 3610
rect 420 3475 435 3595
rect 465 3475 480 3595
rect 420 3460 480 3475
rect 540 3595 600 3610
rect 540 3475 555 3595
rect 585 3475 600 3595
rect 540 3460 600 3475
rect 660 3595 720 3610
rect 660 3475 675 3595
rect 705 3475 720 3595
rect 660 3460 720 3475
rect 780 3595 840 3610
rect 780 3475 795 3595
rect 825 3475 840 3595
rect 780 3460 840 3475
rect 900 3595 960 3610
rect 900 3475 915 3595
rect 945 3475 960 3595
rect 900 3460 960 3475
rect 1020 3595 1080 3610
rect 1020 3475 1035 3595
rect 1065 3475 1080 3595
rect 1020 3460 1080 3475
rect 1140 3595 1200 3610
rect 1140 3475 1155 3595
rect 1185 3475 1200 3595
rect 1140 3460 1200 3475
rect 1260 3595 1320 3610
rect 1260 3475 1275 3595
rect 1305 3475 1320 3595
rect 1260 3460 1320 3475
rect 1380 3595 1440 3610
rect 1380 3475 1395 3595
rect 1425 3475 1440 3595
rect 1380 3460 1440 3475
rect 1500 3595 1560 3610
rect 1500 3475 1515 3595
rect 1545 3475 1560 3595
rect 1500 3460 1560 3475
rect 1620 3595 1680 3610
rect 1620 3475 1635 3595
rect 1665 3475 1680 3595
rect 1620 3460 1680 3475
rect 1740 3595 1800 3610
rect 1740 3475 1755 3595
rect 1785 3475 1800 3595
rect 1740 3460 1800 3475
rect 1860 3595 1920 3610
rect 1860 3475 1875 3595
rect 1905 3475 1920 3595
rect 1860 3460 1920 3475
rect 1980 3595 2040 3610
rect 1980 3475 1995 3595
rect 2025 3475 2040 3595
rect 1980 3460 2040 3475
rect -180 2565 -120 2580
rect -180 2445 -165 2565
rect -135 2445 -120 2565
rect -180 2430 -120 2445
rect -60 2565 0 2580
rect -60 2445 -45 2565
rect -15 2445 0 2565
rect -60 2430 0 2445
rect 60 2565 120 2580
rect 60 2445 75 2565
rect 105 2445 120 2565
rect 60 2430 120 2445
rect 180 2565 240 2580
rect 180 2445 195 2565
rect 225 2445 240 2565
rect 180 2430 240 2445
rect 300 2565 360 2580
rect 300 2445 315 2565
rect 345 2445 360 2565
rect 300 2430 360 2445
rect 420 2565 480 2580
rect 420 2445 435 2565
rect 465 2445 480 2565
rect 420 2430 480 2445
rect 540 2565 600 2580
rect 540 2445 555 2565
rect 585 2445 600 2565
rect 540 2430 600 2445
rect 660 2565 720 2580
rect 660 2445 675 2565
rect 705 2445 720 2565
rect 660 2430 720 2445
rect 780 2565 840 2580
rect 780 2445 795 2565
rect 825 2445 840 2565
rect 780 2430 840 2445
rect 900 2565 960 2580
rect 900 2445 915 2565
rect 945 2445 960 2565
rect 900 2430 960 2445
rect 1020 2565 1080 2580
rect 1020 2445 1035 2565
rect 1065 2445 1080 2565
rect 1020 2430 1080 2445
rect 1140 2565 1200 2580
rect 1140 2445 1155 2565
rect 1185 2445 1200 2565
rect 1140 2430 1200 2445
rect 1260 2565 1320 2580
rect 1260 2445 1275 2565
rect 1305 2445 1320 2565
rect 1260 2430 1320 2445
rect 1380 2565 1440 2580
rect 1380 2445 1395 2565
rect 1425 2445 1440 2565
rect 1380 2430 1440 2445
rect 1500 2565 1560 2580
rect 1500 2445 1515 2565
rect 1545 2445 1560 2565
rect 1500 2430 1560 2445
rect 1620 2565 1680 2580
rect 1620 2445 1635 2565
rect 1665 2445 1680 2565
rect 1620 2430 1680 2445
rect 1740 2565 1800 2580
rect 1740 2445 1755 2565
rect 1785 2445 1800 2565
rect 1740 2430 1800 2445
rect 1860 2565 1920 2580
rect 1860 2445 1875 2565
rect 1905 2445 1920 2565
rect 1860 2430 1920 2445
rect 1980 2565 2040 2580
rect 1980 2445 1995 2565
rect 2025 2445 2040 2565
rect 1980 2430 2040 2445
<< pdiff >>
rect -180 4760 -120 4775
rect -180 4640 -165 4760
rect -135 4640 -120 4760
rect -180 4625 -120 4640
rect -60 4760 0 4775
rect -60 4640 -45 4760
rect -15 4640 0 4760
rect -60 4625 0 4640
rect 60 4760 120 4775
rect 60 4640 75 4760
rect 105 4640 120 4760
rect 60 4625 120 4640
rect 180 4760 240 4775
rect 180 4640 195 4760
rect 225 4640 240 4760
rect 180 4625 240 4640
rect 300 4760 360 4775
rect 300 4640 315 4760
rect 345 4640 360 4760
rect 300 4625 360 4640
rect 420 4760 480 4775
rect 420 4640 435 4760
rect 465 4640 480 4760
rect 420 4625 480 4640
rect 540 4760 600 4775
rect 540 4640 555 4760
rect 585 4640 600 4760
rect 540 4625 600 4640
rect 660 4760 720 4775
rect 660 4640 675 4760
rect 705 4640 720 4760
rect 660 4625 720 4640
rect 780 4760 840 4775
rect 780 4640 795 4760
rect 825 4640 840 4760
rect 780 4625 840 4640
rect 900 4760 960 4775
rect 900 4640 915 4760
rect 945 4640 960 4760
rect 900 4625 960 4640
rect 1020 4760 1080 4775
rect 1020 4640 1035 4760
rect 1065 4640 1080 4760
rect 1020 4625 1080 4640
rect 1140 4760 1200 4775
rect 1140 4640 1155 4760
rect 1185 4640 1200 4760
rect 1140 4625 1200 4640
rect 1260 4760 1320 4775
rect 1260 4640 1275 4760
rect 1305 4640 1320 4760
rect 1260 4625 1320 4640
rect 1380 4760 1440 4775
rect 1380 4640 1395 4760
rect 1425 4640 1440 4760
rect 1380 4625 1440 4640
rect 1500 4760 1560 4775
rect 1500 4640 1515 4760
rect 1545 4640 1560 4760
rect 1500 4625 1560 4640
rect 1620 4760 1680 4775
rect 1620 4640 1635 4760
rect 1665 4640 1680 4760
rect 1620 4625 1680 4640
rect 1740 4760 1800 4775
rect 1740 4640 1755 4760
rect 1785 4640 1800 4760
rect 1740 4625 1800 4640
rect 1860 4760 1920 4775
rect 1860 4640 1875 4760
rect 1905 4640 1920 4760
rect 1860 4625 1920 4640
rect 1980 4760 2040 4775
rect 1980 4640 1995 4760
rect 2025 4640 2040 4760
rect 1980 4625 2040 4640
rect -180 4035 -120 4050
rect -180 3915 -165 4035
rect -135 3915 -120 4035
rect -180 3900 -120 3915
rect -60 4035 0 4050
rect -60 3915 -45 4035
rect -15 3915 0 4035
rect -60 3900 0 3915
rect 60 4035 120 4050
rect 60 3915 75 4035
rect 105 3915 120 4035
rect 60 3900 120 3915
rect 180 4035 240 4050
rect 180 3915 195 4035
rect 225 3915 240 4035
rect 180 3900 240 3915
rect 300 4035 360 4050
rect 300 3915 315 4035
rect 345 3915 360 4035
rect 300 3900 360 3915
rect 420 4035 480 4050
rect 420 3915 435 4035
rect 465 3915 480 4035
rect 420 3900 480 3915
rect 540 4035 600 4050
rect 540 3915 555 4035
rect 585 3915 600 4035
rect 540 3900 600 3915
rect 660 4035 720 4050
rect 660 3915 675 4035
rect 705 3915 720 4035
rect 660 3900 720 3915
rect 780 4035 840 4050
rect 780 3915 795 4035
rect 825 3915 840 4035
rect 780 3900 840 3915
rect 900 4035 960 4050
rect 900 3915 915 4035
rect 945 3915 960 4035
rect 900 3900 960 3915
rect 1020 4035 1080 4050
rect 1020 3915 1035 4035
rect 1065 3915 1080 4035
rect 1020 3900 1080 3915
rect 1140 4035 1200 4050
rect 1140 3915 1155 4035
rect 1185 3915 1200 4035
rect 1140 3900 1200 3915
rect 1260 4035 1320 4050
rect 1260 3915 1275 4035
rect 1305 3915 1320 4035
rect 1260 3900 1320 3915
rect 1380 4035 1440 4050
rect 1380 3915 1395 4035
rect 1425 3915 1440 4035
rect 1380 3900 1440 3915
rect 1500 4035 1560 4050
rect 1500 3915 1515 4035
rect 1545 3915 1560 4035
rect 1500 3900 1560 3915
rect 1620 4035 1680 4050
rect 1620 3915 1635 4035
rect 1665 3915 1680 4035
rect 1620 3900 1680 3915
rect 1740 4035 1800 4050
rect 1740 3915 1755 4035
rect 1785 3915 1800 4035
rect 1740 3900 1800 3915
rect 1860 4035 1920 4050
rect 1860 3915 1875 4035
rect 1905 3915 1920 4035
rect 1860 3900 1920 3915
rect 1980 4035 2040 4050
rect 1980 3915 1995 4035
rect 2025 3915 2040 4035
rect 1980 3900 2040 3915
rect -180 3100 -120 3115
rect -180 2980 -165 3100
rect -135 2980 -120 3100
rect -180 2965 -120 2980
rect -60 3100 0 3115
rect -60 2980 -45 3100
rect -15 2980 0 3100
rect -60 2965 0 2980
rect 60 3100 120 3115
rect 60 2980 75 3100
rect 105 2980 120 3100
rect 60 2965 120 2980
rect 180 3100 240 3115
rect 180 2980 195 3100
rect 225 2980 240 3100
rect 180 2965 240 2980
rect 300 3100 360 3115
rect 300 2980 315 3100
rect 345 2980 360 3100
rect 300 2965 360 2980
rect 420 3100 480 3115
rect 420 2980 435 3100
rect 465 2980 480 3100
rect 420 2965 480 2980
rect 540 3100 600 3115
rect 540 2980 555 3100
rect 585 2980 600 3100
rect 540 2965 600 2980
rect 660 3100 720 3115
rect 660 2980 675 3100
rect 705 2980 720 3100
rect 660 2965 720 2980
rect 780 3100 840 3115
rect 780 2980 795 3100
rect 825 2980 840 3100
rect 780 2965 840 2980
rect 900 3100 960 3115
rect 900 2980 915 3100
rect 945 2980 960 3100
rect 900 2965 960 2980
rect 1020 3100 1080 3115
rect 1020 2980 1035 3100
rect 1065 2980 1080 3100
rect 1020 2965 1080 2980
rect 1140 3100 1200 3115
rect 1140 2980 1155 3100
rect 1185 2980 1200 3100
rect 1140 2965 1200 2980
rect 1260 3100 1320 3115
rect 1260 2980 1275 3100
rect 1305 2980 1320 3100
rect 1260 2965 1320 2980
rect 1380 3100 1440 3115
rect 1380 2980 1395 3100
rect 1425 2980 1440 3100
rect 1380 2965 1440 2980
rect 1500 3100 1560 3115
rect 1500 2980 1515 3100
rect 1545 2980 1560 3100
rect 1500 2965 1560 2980
rect 1620 3100 1680 3115
rect 1620 2980 1635 3100
rect 1665 2980 1680 3100
rect 1620 2965 1680 2980
rect 1740 3100 1800 3115
rect 1740 2980 1755 3100
rect 1785 2980 1800 3100
rect 1740 2965 1800 2980
rect 1860 3100 1920 3115
rect 1860 2980 1875 3100
rect 1905 2980 1920 3100
rect 1860 2965 1920 2980
rect 1980 3100 2040 3115
rect 1980 2980 1995 3100
rect 2025 2980 2040 3100
rect 1980 2965 2040 2980
<< ndiffc >>
rect -165 4310 -135 4430
rect -45 4310 -15 4430
rect 75 4310 105 4430
rect 195 4310 225 4430
rect 315 4310 345 4430
rect 435 4310 465 4430
rect 555 4310 585 4430
rect 675 4310 705 4430
rect 795 4310 825 4430
rect 915 4310 945 4430
rect 1035 4310 1065 4430
rect 1155 4310 1185 4430
rect 1275 4310 1305 4430
rect 1395 4310 1425 4430
rect 1515 4310 1545 4430
rect 1635 4310 1665 4430
rect 1755 4310 1785 4430
rect 1875 4310 1905 4430
rect 1995 4310 2025 4430
rect -165 3475 -135 3595
rect -45 3475 -15 3595
rect 75 3475 105 3595
rect 195 3475 225 3595
rect 315 3475 345 3595
rect 435 3475 465 3595
rect 555 3475 585 3595
rect 675 3475 705 3595
rect 795 3475 825 3595
rect 915 3475 945 3595
rect 1035 3475 1065 3595
rect 1155 3475 1185 3595
rect 1275 3475 1305 3595
rect 1395 3475 1425 3595
rect 1515 3475 1545 3595
rect 1635 3475 1665 3595
rect 1755 3475 1785 3595
rect 1875 3475 1905 3595
rect 1995 3475 2025 3595
rect -165 2445 -135 2565
rect -45 2445 -15 2565
rect 75 2445 105 2565
rect 195 2445 225 2565
rect 315 2445 345 2565
rect 435 2445 465 2565
rect 555 2445 585 2565
rect 675 2445 705 2565
rect 795 2445 825 2565
rect 915 2445 945 2565
rect 1035 2445 1065 2565
rect 1155 2445 1185 2565
rect 1275 2445 1305 2565
rect 1395 2445 1425 2565
rect 1515 2445 1545 2565
rect 1635 2445 1665 2565
rect 1755 2445 1785 2565
rect 1875 2445 1905 2565
rect 1995 2445 2025 2565
<< pdiffc >>
rect -165 4640 -135 4760
rect -45 4640 -15 4760
rect 75 4640 105 4760
rect 195 4640 225 4760
rect 315 4640 345 4760
rect 435 4640 465 4760
rect 555 4640 585 4760
rect 675 4640 705 4760
rect 795 4640 825 4760
rect 915 4640 945 4760
rect 1035 4640 1065 4760
rect 1155 4640 1185 4760
rect 1275 4640 1305 4760
rect 1395 4640 1425 4760
rect 1515 4640 1545 4760
rect 1635 4640 1665 4760
rect 1755 4640 1785 4760
rect 1875 4640 1905 4760
rect 1995 4640 2025 4760
rect -165 3915 -135 4035
rect -45 3915 -15 4035
rect 75 3915 105 4035
rect 195 3915 225 4035
rect 315 3915 345 4035
rect 435 3915 465 4035
rect 555 3915 585 4035
rect 675 3915 705 4035
rect 795 3915 825 4035
rect 915 3915 945 4035
rect 1035 3915 1065 4035
rect 1155 3915 1185 4035
rect 1275 3915 1305 4035
rect 1395 3915 1425 4035
rect 1515 3915 1545 4035
rect 1635 3915 1665 4035
rect 1755 3915 1785 4035
rect 1875 3915 1905 4035
rect 1995 3915 2025 4035
rect -165 2980 -135 3100
rect -45 2980 -15 3100
rect 75 2980 105 3100
rect 195 2980 225 3100
rect 315 2980 345 3100
rect 435 2980 465 3100
rect 555 2980 585 3100
rect 675 2980 705 3100
rect 795 2980 825 3100
rect 915 2980 945 3100
rect 1035 2980 1065 3100
rect 1155 2980 1185 3100
rect 1275 2980 1305 3100
rect 1395 2980 1425 3100
rect 1515 2980 1545 3100
rect 1635 2980 1665 3100
rect 1755 2980 1785 3100
rect 1875 2980 1905 3100
rect 1995 2980 2025 3100
<< psubdiff >>
rect 165 4525 225 4540
rect 165 4495 180 4525
rect 210 4495 225 4525
rect 165 4480 225 4495
rect 1720 4540 1780 4555
rect 1720 4510 1735 4540
rect 1765 4510 1780 4540
rect 1720 4495 1780 4510
rect 165 3755 225 3770
rect 165 3720 180 3755
rect 210 3720 225 3755
rect 1675 3745 1735 3760
rect 165 3705 225 3720
rect 1675 3710 1690 3745
rect 1720 3710 1735 3745
rect 1675 3695 1735 3710
rect 455 2730 575 2745
rect 455 2640 470 2730
rect 560 2640 575 2730
rect 1300 2730 1420 2745
rect 455 2625 575 2640
rect 1300 2640 1315 2730
rect 1405 2640 1420 2730
rect 1300 2625 1420 2640
<< nsubdiff >>
rect 350 4540 410 4560
rect 350 4515 365 4540
rect 395 4515 410 4540
rect 350 4500 410 4515
rect 1530 4545 1590 4560
rect 1530 4525 1550 4545
rect 1570 4525 1590 4545
rect 1530 4510 1590 4525
rect 360 3835 420 3850
rect 360 3800 375 3835
rect 405 3800 420 3835
rect 1440 3825 1500 3840
rect 360 3785 420 3800
rect 1440 3790 1455 3825
rect 1485 3790 1500 3825
rect 1440 3775 1500 3790
rect 235 2870 355 2885
rect 235 2780 250 2870
rect 340 2780 355 2870
rect 1625 2870 1745 2885
rect 235 2765 355 2780
rect 1625 2780 1640 2870
rect 1730 2780 1745 2870
rect 1625 2765 1745 2780
<< psubdiffcont >>
rect 180 4495 210 4525
rect 1735 4510 1765 4540
rect 180 3720 210 3755
rect 1690 3710 1720 3745
rect 470 2640 560 2730
rect 1315 2640 1405 2730
<< nsubdiffcont >>
rect 365 4515 395 4540
rect 1550 4525 1570 4545
rect 375 3800 405 3835
rect 1455 3790 1485 3825
rect 250 2780 340 2870
rect 1640 2780 1730 2870
<< poly >>
rect -240 4815 1380 4830
rect -120 4775 -60 4790
rect 0 4775 60 4790
rect 120 4775 180 4790
rect 240 4775 300 4790
rect 360 4775 420 4790
rect 480 4775 540 4815
rect 600 4775 660 4790
rect 720 4775 780 4790
rect 840 4775 900 4790
rect 960 4775 1020 4790
rect 1080 4775 1140 4790
rect 1200 4775 1260 4790
rect 1320 4775 1380 4815
rect 1440 4775 1500 4790
rect 1560 4775 1620 4790
rect 1680 4775 1740 4790
rect 1800 4775 1860 4790
rect 1920 4775 1980 4790
rect -120 4610 -60 4625
rect 0 4610 60 4625
rect 120 4610 180 4625
rect 240 4610 300 4625
rect 360 4610 420 4625
rect -175 4600 420 4610
rect -175 4580 -165 4600
rect -70 4580 -45 4600
rect 50 4580 75 4600
rect 170 4580 195 4600
rect 290 4580 315 4600
rect 410 4580 420 4600
rect -175 4570 420 4580
rect -120 4445 -60 4460
rect 0 4445 60 4460
rect 120 4445 180 4460
rect 240 4445 300 4460
rect 360 4445 420 4460
rect 480 4445 540 4625
rect 600 4610 660 4625
rect 720 4585 780 4625
rect 600 4570 780 4585
rect 600 4445 660 4570
rect 840 4540 900 4625
rect 960 4540 1020 4625
rect 1080 4585 1140 4625
rect 1200 4610 1260 4625
rect 1080 4570 1260 4585
rect 840 4530 1020 4540
rect 840 4525 920 4530
rect 910 4510 920 4525
rect 940 4525 1020 4530
rect 940 4510 950 4525
rect 910 4500 950 4510
rect 720 4445 780 4460
rect 840 4445 900 4460
rect 960 4445 1020 4460
rect 1080 4445 1140 4460
rect 1200 4445 1260 4570
rect 1320 4445 1380 4625
rect 1440 4610 1500 4625
rect 1560 4610 1620 4625
rect 1680 4610 1740 4625
rect 1800 4610 1860 4625
rect 1920 4610 1980 4625
rect 1440 4600 2035 4610
rect 1440 4580 1450 4600
rect 1545 4580 1570 4600
rect 1665 4580 1690 4600
rect 1785 4580 1810 4600
rect 1905 4580 1930 4600
rect 2025 4580 2035 4600
rect 1440 4570 2035 4580
rect 2020 4490 2060 4500
rect 2020 4470 2030 4490
rect 2050 4475 2060 4490
rect 2050 4470 2075 4475
rect 2020 4460 2075 4470
rect 1440 4445 1500 4460
rect 1560 4445 1620 4460
rect 1680 4445 1740 4460
rect 1800 4445 1860 4460
rect 1920 4445 1980 4460
rect -120 4280 -60 4295
rect 0 4280 60 4295
rect 120 4280 180 4295
rect 240 4280 300 4295
rect 360 4280 420 4295
rect 480 4280 540 4295
rect -175 4270 420 4280
rect -175 4250 -165 4270
rect -70 4250 -45 4270
rect 50 4250 75 4270
rect 170 4250 195 4270
rect 290 4250 315 4270
rect 410 4250 420 4270
rect -175 4240 420 4250
rect 600 4205 660 4295
rect 720 4280 780 4295
rect -240 4190 660 4205
rect 840 4255 900 4295
rect 960 4255 1020 4295
rect 1080 4280 1140 4295
rect 1200 4280 1260 4295
rect 1320 4280 1380 4295
rect 1440 4280 1500 4295
rect 1560 4280 1620 4295
rect 1680 4280 1740 4295
rect 1800 4280 1860 4295
rect 1920 4280 1980 4295
rect 840 4240 1020 4255
rect 1440 4270 2035 4280
rect 1440 4250 1450 4270
rect 1545 4250 1570 4270
rect 1665 4250 1690 4270
rect 1785 4250 1810 4270
rect 1905 4250 1930 4270
rect 2025 4250 2035 4270
rect 1440 4240 2035 4250
rect 840 4165 855 4240
rect -220 4150 855 4165
rect -220 3690 -205 4150
rect 2060 4105 2075 4460
rect 360 4090 2075 4105
rect -120 4050 -60 4065
rect 0 4050 60 4065
rect 120 4050 180 4065
rect 240 4050 300 4065
rect 360 4050 420 4090
rect 480 4050 540 4065
rect 600 4050 660 4065
rect 720 4050 780 4090
rect 840 4050 900 4065
rect 960 4050 1020 4065
rect 1080 4050 1140 4090
rect 1200 4050 1260 4065
rect 1320 4050 1380 4065
rect 1440 4050 1500 4090
rect 1560 4050 1620 4065
rect 1680 4050 1740 4065
rect 1800 4050 1860 4065
rect 1920 4050 1980 4065
rect -120 3885 -60 3900
rect 0 3885 60 3900
rect 120 3885 180 3900
rect 240 3885 300 3900
rect 360 3885 420 3900
rect -175 3875 300 3885
rect -175 3855 -165 3875
rect -70 3855 -45 3875
rect 50 3855 75 3875
rect 170 3855 195 3875
rect 290 3855 300 3875
rect -175 3845 300 3855
rect 480 3875 540 3900
rect 600 3885 660 3900
rect 720 3885 780 3900
rect 480 3855 490 3875
rect 530 3855 540 3875
rect 480 3845 540 3855
rect 840 3875 900 3900
rect 840 3855 850 3875
rect 890 3855 900 3875
rect 840 3845 900 3855
rect 960 3875 1020 3900
rect 1080 3885 1140 3900
rect 1200 3885 1260 3900
rect 960 3855 970 3875
rect 1010 3855 1020 3875
rect 960 3845 1020 3855
rect 1320 3875 1380 3900
rect 1440 3885 1500 3900
rect 1560 3885 1620 3900
rect 1680 3885 1740 3900
rect 1800 3885 1860 3900
rect 1920 3885 1980 3900
rect 1320 3855 1330 3875
rect 1370 3855 1380 3875
rect 1320 3845 1380 3855
rect 1560 3875 2035 3885
rect 1560 3855 1570 3875
rect 1665 3855 1690 3875
rect 1785 3855 1810 3875
rect 1905 3855 1930 3875
rect 2025 3855 2035 3875
rect 1560 3845 2035 3855
rect 910 3815 950 3825
rect 910 3795 920 3815
rect 940 3795 950 3815
rect 910 3785 950 3795
rect 920 3725 940 3785
rect 910 3715 950 3725
rect 910 3695 920 3715
rect 940 3695 950 3715
rect -220 3675 420 3690
rect 910 3685 950 3695
rect -120 3610 -60 3625
rect 0 3610 60 3625
rect 120 3610 180 3625
rect 240 3610 300 3625
rect 360 3610 420 3675
rect 480 3655 540 3665
rect 480 3635 490 3655
rect 530 3635 540 3655
rect 480 3610 540 3635
rect 840 3655 900 3665
rect 840 3635 850 3655
rect 890 3635 900 3655
rect 600 3610 660 3625
rect 720 3610 780 3625
rect 840 3610 900 3635
rect 960 3655 1020 3665
rect 960 3635 970 3655
rect 1010 3635 1020 3655
rect 960 3610 1020 3635
rect 1320 3655 1380 3665
rect 1320 3635 1330 3655
rect 1370 3635 1380 3655
rect 1080 3610 1140 3625
rect 1200 3610 1260 3625
rect 1320 3610 1380 3635
rect 1440 3610 1500 3625
rect 1560 3610 1620 3625
rect 1680 3610 1740 3625
rect 1800 3610 1860 3625
rect 1920 3610 1980 3625
rect -120 3445 -60 3460
rect 0 3445 60 3460
rect 120 3445 180 3460
rect 240 3445 300 3460
rect -175 3435 300 3445
rect -175 3415 -165 3435
rect -70 3415 -45 3435
rect 50 3415 75 3435
rect 170 3415 195 3435
rect 290 3415 300 3435
rect -175 3405 300 3415
rect 360 3420 420 3460
rect 480 3445 540 3460
rect 600 3445 660 3460
rect 720 3420 780 3460
rect 840 3445 900 3460
rect 960 3445 1020 3460
rect 1080 3420 1140 3460
rect 1200 3445 1260 3460
rect 1320 3445 1380 3460
rect 1440 3420 1500 3460
rect 360 3405 1500 3420
rect 1560 3445 1620 3460
rect 1680 3445 1740 3460
rect 1800 3445 1860 3460
rect 1920 3445 1980 3460
rect 1560 3435 2035 3445
rect 1560 3415 1570 3435
rect 1665 3415 1690 3435
rect 1785 3415 1810 3435
rect 1905 3415 1930 3435
rect 2025 3415 2035 3435
rect 1560 3405 2035 3415
rect 440 3190 460 3405
rect 430 3180 470 3190
rect 430 3160 440 3180
rect 460 3160 470 3180
rect 2060 3175 2075 4090
rect 430 3150 470 3160
rect 1800 3160 2075 3175
rect -120 3115 -60 3130
rect 0 3115 60 3130
rect 120 3115 180 3130
rect 240 3115 300 3130
rect 360 3115 420 3130
rect 480 3115 540 3130
rect 600 3115 660 3130
rect 720 3115 780 3130
rect 840 3115 900 3130
rect 960 3115 1020 3130
rect 1080 3115 1140 3130
rect 1200 3115 1260 3130
rect 1320 3115 1380 3130
rect 1440 3115 1500 3130
rect 1560 3115 1620 3130
rect 1680 3115 1740 3130
rect 1800 3115 1860 3160
rect 1920 3115 1980 3130
rect -120 2950 -60 2965
rect -175 2940 -60 2950
rect -175 2920 -165 2940
rect -70 2920 -60 2940
rect -175 2910 -60 2920
rect 0 2925 60 2965
rect 120 2925 180 2965
rect 240 2925 300 2965
rect 360 2950 420 2965
rect 480 2925 540 2965
rect 600 2925 660 2965
rect 720 2950 780 2965
rect 840 2925 900 2965
rect 960 2925 1020 2965
rect 1080 2950 1140 2965
rect 1200 2925 1260 2965
rect 1320 2925 1380 2965
rect 1440 2950 1500 2965
rect 1560 2925 1620 2965
rect 1680 2925 1740 2965
rect 1800 2925 1860 2965
rect 0 2910 1860 2925
rect 1920 2950 1980 2965
rect 1920 2940 2035 2950
rect 1920 2920 1930 2940
rect 2025 2920 2035 2940
rect 1920 2910 2035 2920
rect 785 2875 835 2885
rect 785 2850 795 2875
rect 825 2855 835 2875
rect 1025 2875 1075 2885
rect 1025 2855 1035 2875
rect 825 2850 1035 2855
rect 1065 2850 1075 2875
rect 425 2835 475 2850
rect 785 2840 1075 2850
rect 425 2810 435 2835
rect 465 2815 475 2835
rect 1385 2835 1435 2850
rect 1385 2815 1395 2835
rect 465 2810 1395 2815
rect 1425 2810 1435 2835
rect 425 2800 1435 2810
rect 920 2665 940 2800
rect 905 2655 955 2665
rect 905 2630 915 2655
rect 945 2630 955 2655
rect 905 2620 955 2630
rect -120 2580 -60 2595
rect 0 2580 60 2595
rect 120 2580 180 2595
rect 240 2580 300 2595
rect 360 2580 420 2595
rect 480 2580 540 2595
rect 600 2580 660 2595
rect 720 2580 780 2595
rect 840 2580 900 2595
rect 960 2580 1020 2595
rect 1080 2580 1140 2595
rect 1200 2580 1260 2595
rect 1320 2580 1380 2595
rect 1440 2580 1500 2595
rect 1560 2580 1620 2595
rect 1680 2580 1740 2595
rect 1800 2580 1860 2595
rect 1920 2580 1980 2595
rect -120 2415 -60 2430
rect -175 2405 -60 2415
rect -175 2385 -165 2405
rect -70 2385 -60 2405
rect -175 2375 -60 2385
rect 0 2390 60 2430
rect 120 2390 180 2430
rect 240 2390 300 2430
rect 360 2415 420 2430
rect 480 2390 540 2430
rect 600 2390 660 2430
rect 720 2415 780 2430
rect 840 2395 900 2430
rect 960 2395 1020 2430
rect 1080 2415 1140 2430
rect 840 2390 1020 2395
rect 1200 2390 1260 2430
rect 1320 2390 1380 2430
rect 1440 2415 1500 2430
rect 1560 2390 1620 2430
rect 1680 2390 1740 2430
rect 1800 2390 1860 2430
rect 0 2385 1860 2390
rect 0 2375 920 2385
rect 910 2365 920 2375
rect 940 2375 1860 2385
rect 1920 2415 1980 2430
rect 1920 2405 2035 2415
rect 1920 2385 1930 2405
rect 2025 2385 2035 2405
rect 1920 2375 2035 2385
rect 940 2365 950 2375
rect 910 2355 950 2365
<< polycont >>
rect -165 4580 -70 4600
rect -45 4580 50 4600
rect 75 4580 170 4600
rect 195 4580 290 4600
rect 315 4580 410 4600
rect 920 4510 940 4530
rect 1450 4580 1545 4600
rect 1570 4580 1665 4600
rect 1690 4580 1785 4600
rect 1810 4580 1905 4600
rect 1930 4580 2025 4600
rect 2030 4470 2050 4490
rect -165 4250 -70 4270
rect -45 4250 50 4270
rect 75 4250 170 4270
rect 195 4250 290 4270
rect 315 4250 410 4270
rect 1450 4250 1545 4270
rect 1570 4250 1665 4270
rect 1690 4250 1785 4270
rect 1810 4250 1905 4270
rect 1930 4250 2025 4270
rect -165 3855 -70 3875
rect -45 3855 50 3875
rect 75 3855 170 3875
rect 195 3855 290 3875
rect 490 3855 530 3875
rect 850 3855 890 3875
rect 970 3855 1010 3875
rect 1330 3855 1370 3875
rect 1570 3855 1665 3875
rect 1690 3855 1785 3875
rect 1810 3855 1905 3875
rect 1930 3855 2025 3875
rect 920 3795 940 3815
rect 920 3695 940 3715
rect 490 3635 530 3655
rect 850 3635 890 3655
rect 970 3635 1010 3655
rect 1330 3635 1370 3655
rect -165 3415 -70 3435
rect -45 3415 50 3435
rect 75 3415 170 3435
rect 195 3415 290 3435
rect 1570 3415 1665 3435
rect 1690 3415 1785 3435
rect 1810 3415 1905 3435
rect 1930 3415 2025 3435
rect 440 3160 460 3180
rect -165 2920 -70 2940
rect 1930 2920 2025 2940
rect 795 2850 825 2875
rect 1035 2850 1065 2875
rect 435 2810 465 2835
rect 1395 2810 1425 2835
rect 915 2630 945 2655
rect -165 2385 -70 2405
rect 920 2365 940 2385
rect 1930 2385 2025 2405
<< locali >>
rect 425 4850 1435 4870
rect 425 4815 475 4850
rect -225 4795 475 4815
rect -225 3330 -205 4795
rect -175 4760 -125 4770
rect -175 4640 -165 4760
rect -135 4640 -125 4760
rect -175 4610 -125 4640
rect -55 4760 -5 4770
rect -55 4640 -45 4760
rect -15 4640 -5 4760
rect -55 4610 -5 4640
rect 65 4760 115 4770
rect 65 4640 75 4760
rect 105 4640 115 4760
rect 65 4610 115 4640
rect 185 4760 235 4770
rect 185 4640 195 4760
rect 225 4640 235 4760
rect 185 4610 235 4640
rect 305 4760 355 4770
rect 305 4640 315 4760
rect 345 4640 355 4760
rect 305 4610 355 4640
rect 425 4760 475 4795
rect 425 4640 435 4760
rect 465 4640 475 4760
rect 425 4630 475 4640
rect 545 4810 1315 4830
rect 545 4760 595 4810
rect 545 4640 555 4760
rect 585 4640 595 4760
rect 545 4630 595 4640
rect 665 4760 715 4770
rect 665 4640 675 4760
rect 705 4640 715 4760
rect -175 4600 420 4610
rect -175 4580 -165 4600
rect -70 4580 -45 4600
rect 50 4580 75 4600
rect 170 4580 195 4600
rect 290 4580 315 4600
rect 410 4580 420 4600
rect -175 4570 420 4580
rect 665 4585 715 4640
rect 785 4760 835 4810
rect 785 4640 795 4760
rect 825 4640 835 4760
rect 785 4630 835 4640
rect 905 4760 955 4770
rect 905 4640 915 4760
rect 945 4640 955 4760
rect 905 4630 955 4640
rect 1025 4760 1075 4810
rect 1025 4640 1035 4760
rect 1065 4640 1075 4760
rect 1025 4630 1075 4640
rect 1145 4760 1195 4770
rect 1145 4640 1155 4760
rect 1185 4640 1195 4760
rect 1145 4585 1195 4640
rect 1265 4760 1315 4810
rect 1265 4640 1275 4760
rect 1305 4640 1315 4760
rect 1265 4630 1315 4640
rect 1385 4760 1435 4850
rect 1385 4640 1395 4760
rect 1425 4640 1435 4760
rect 1385 4630 1435 4640
rect 1505 4760 1555 4770
rect 1505 4640 1515 4760
rect 1545 4640 1555 4760
rect 1505 4610 1555 4640
rect 1625 4760 1675 4770
rect 1625 4640 1635 4760
rect 1665 4640 1675 4760
rect 1625 4610 1675 4640
rect 1745 4760 1795 4770
rect 1745 4640 1755 4760
rect 1785 4640 1795 4760
rect 1745 4610 1795 4640
rect 1865 4760 1915 4770
rect 1865 4640 1875 4760
rect 1905 4640 1915 4760
rect 1865 4610 1915 4640
rect 1985 4760 2035 4770
rect 1985 4640 1995 4760
rect 2025 4640 2035 4760
rect 1985 4610 2035 4640
rect 665 4565 1195 4585
rect 1440 4600 2035 4610
rect 1440 4580 1450 4600
rect 1545 4580 1570 4600
rect 1665 4580 1690 4600
rect 1785 4580 1810 4600
rect 1905 4580 1930 4600
rect 2025 4580 2035 4600
rect 1440 4570 2035 4580
rect 355 4540 405 4550
rect 1540 4545 1580 4550
rect 170 4525 220 4535
rect 170 4495 180 4525
rect 210 4495 220 4525
rect 355 4515 365 4540
rect 395 4515 405 4540
rect 355 4505 405 4515
rect 910 4530 950 4540
rect 910 4510 920 4530
rect 940 4520 950 4530
rect 1540 4525 1550 4545
rect 1570 4525 1580 4545
rect 1540 4520 1580 4525
rect 1725 4540 1775 4550
rect 940 4510 1235 4520
rect 910 4500 1235 4510
rect 1725 4510 1735 4540
rect 1765 4510 1775 4540
rect 1725 4500 1775 4510
rect 170 4485 220 4495
rect 1215 4480 1235 4500
rect 2020 4490 2060 4500
rect 2020 4480 2030 4490
rect 665 4460 1195 4480
rect 1215 4470 2030 4480
rect 2050 4470 2060 4490
rect 1215 4460 2060 4470
rect -175 4430 -125 4440
rect -175 4310 -165 4430
rect -135 4310 -125 4430
rect -175 4280 -125 4310
rect -55 4430 -5 4440
rect -55 4310 -45 4430
rect -15 4310 -5 4430
rect -55 4280 -5 4310
rect 65 4430 115 4440
rect 65 4310 75 4430
rect 105 4310 115 4430
rect 65 4280 115 4310
rect 185 4430 235 4440
rect 185 4310 195 4430
rect 225 4310 235 4430
rect 185 4280 235 4310
rect 305 4430 355 4440
rect 305 4310 315 4430
rect 345 4310 355 4430
rect 305 4280 355 4310
rect 425 4430 475 4440
rect 425 4310 435 4430
rect 465 4310 475 4430
rect 425 4300 475 4310
rect -175 4270 420 4280
rect -175 4250 -165 4270
rect -70 4250 -45 4270
rect 50 4250 75 4270
rect 170 4250 195 4270
rect 290 4250 315 4270
rect 410 4250 420 4270
rect -175 4240 420 4250
rect 455 4235 475 4300
rect 545 4430 595 4440
rect 545 4310 555 4430
rect 585 4310 595 4430
rect 545 4275 595 4310
rect 665 4430 715 4460
rect 665 4310 675 4430
rect 705 4310 715 4430
rect 665 4300 715 4310
rect 785 4430 835 4440
rect 785 4310 795 4430
rect 825 4310 835 4430
rect 785 4275 835 4310
rect 905 4430 955 4440
rect 905 4310 915 4430
rect 945 4310 955 4430
rect 905 4300 955 4310
rect 1025 4430 1075 4440
rect 1025 4310 1035 4430
rect 1065 4310 1075 4430
rect 1025 4275 1075 4310
rect 1145 4430 1195 4460
rect 1145 4310 1155 4430
rect 1185 4310 1195 4430
rect 1145 4300 1195 4310
rect 1265 4430 1315 4440
rect 1265 4310 1275 4430
rect 1305 4310 1315 4430
rect 1265 4275 1315 4310
rect 545 4255 1315 4275
rect 1385 4430 1435 4440
rect 1385 4310 1395 4430
rect 1425 4310 1435 4430
rect 1385 4300 1435 4310
rect 1505 4430 1555 4440
rect 1505 4310 1515 4430
rect 1545 4310 1555 4430
rect 1385 4235 1405 4300
rect 1505 4280 1555 4310
rect 1625 4430 1675 4440
rect 1625 4310 1635 4430
rect 1665 4310 1675 4430
rect 1625 4280 1675 4310
rect 1745 4430 1795 4440
rect 1745 4310 1755 4430
rect 1785 4310 1795 4430
rect 1745 4280 1795 4310
rect 1865 4430 1915 4440
rect 1865 4310 1875 4430
rect 1905 4310 1915 4430
rect 1865 4280 1915 4310
rect 1985 4430 2035 4440
rect 1985 4310 1995 4430
rect 2025 4310 2035 4430
rect 1985 4280 2035 4310
rect 1440 4270 2035 4280
rect 1440 4250 1450 4270
rect 1545 4250 1570 4270
rect 1665 4250 1690 4270
rect 1785 4250 1810 4270
rect 1905 4250 1930 4270
rect 2025 4250 2035 4270
rect 1440 4240 2035 4250
rect 455 4215 1405 4235
rect 455 4195 475 4215
rect 1385 4195 1405 4215
rect 455 4175 2080 4195
rect 455 4050 475 4175
rect -175 4035 -125 4045
rect -175 3915 -165 4035
rect -135 3915 -125 4035
rect -175 3885 -125 3915
rect -55 4035 -5 4045
rect -55 3915 -45 4035
rect -15 3915 -5 4035
rect -55 3885 -5 3915
rect 65 4035 115 4045
rect 65 3915 75 4035
rect 105 3915 115 4035
rect 65 3885 115 3915
rect 185 4035 235 4045
rect 185 3915 195 4035
rect 225 3915 235 4035
rect 185 3885 235 3915
rect 305 4035 355 4045
rect 305 3915 315 4035
rect 345 3915 355 4035
rect 305 3905 355 3915
rect 425 4035 475 4050
rect 785 4135 1075 4155
rect 425 3915 435 4035
rect 465 3915 475 4035
rect 425 3905 475 3915
rect 545 4035 595 4045
rect 545 3915 555 4035
rect 585 3915 595 4035
rect 545 3885 595 3915
rect 665 4035 715 4045
rect 665 3915 675 4035
rect 705 3915 715 4035
rect 665 3905 715 3915
rect 785 4035 835 4135
rect 785 3915 795 4035
rect 825 3915 835 4035
rect 785 3905 835 3915
rect 905 4035 955 4045
rect 905 3915 915 4035
rect 945 3915 955 4035
rect 905 3905 955 3915
rect 1025 4035 1075 4135
rect 1385 4050 1405 4175
rect 1025 3915 1035 4035
rect 1065 3915 1075 4035
rect 1025 3905 1075 3915
rect 1145 4035 1195 4045
rect 1145 3915 1155 4035
rect 1185 3915 1195 4035
rect 1145 3905 1195 3915
rect 1265 4035 1315 4045
rect 1265 3915 1275 4035
rect 1305 3915 1315 4035
rect -175 3875 300 3885
rect -175 3855 -165 3875
rect -70 3855 -45 3875
rect 50 3855 75 3875
rect 170 3855 195 3875
rect 290 3855 300 3875
rect -175 3845 300 3855
rect 480 3875 595 3885
rect 480 3855 490 3875
rect 530 3855 595 3875
rect 480 3845 595 3855
rect 840 3875 900 3885
rect 840 3855 850 3875
rect 890 3855 900 3875
rect 840 3845 900 3855
rect 365 3835 415 3845
rect 365 3800 375 3835
rect 405 3800 415 3835
rect 365 3790 415 3800
rect 480 3765 540 3845
rect 840 3765 890 3845
rect 920 3825 940 3905
rect 1265 3885 1315 3915
rect 1385 4035 1435 4050
rect 1385 3915 1395 4035
rect 1425 3915 1435 4035
rect 1385 3905 1435 3915
rect 1505 4035 1555 4045
rect 1505 3915 1515 4035
rect 1545 3915 1555 4035
rect 1505 3905 1555 3915
rect 1625 4035 1675 4045
rect 1625 3915 1635 4035
rect 1665 3915 1675 4035
rect 1625 3885 1675 3915
rect 1745 4035 1795 4045
rect 1745 3915 1755 4035
rect 1785 3915 1795 4035
rect 1745 3885 1795 3915
rect 1865 4035 1915 4045
rect 1865 3915 1875 4035
rect 1905 3915 1915 4035
rect 1865 3885 1915 3915
rect 1985 4035 2035 4045
rect 1985 3915 1995 4035
rect 2025 3915 2035 4035
rect 1985 3885 2035 3915
rect 960 3875 1020 3885
rect 960 3855 970 3875
rect 1010 3855 1020 3875
rect 960 3845 1020 3855
rect 1265 3875 1380 3885
rect 1265 3855 1330 3875
rect 1370 3855 1380 3875
rect 1265 3845 1380 3855
rect 1560 3875 2035 3885
rect 1560 3855 1570 3875
rect 1665 3855 1690 3875
rect 1785 3855 1810 3875
rect 1905 3855 1930 3875
rect 2025 3855 2035 3875
rect 1560 3845 2035 3855
rect 910 3815 950 3825
rect 910 3795 920 3815
rect 940 3795 950 3815
rect 910 3785 950 3795
rect 970 3765 1020 3845
rect 1320 3765 1380 3845
rect 1445 3825 1495 3835
rect 1445 3790 1455 3825
rect 1485 3790 1495 3825
rect 1445 3780 1495 3790
rect 170 3755 220 3765
rect 170 3720 180 3755
rect 210 3720 220 3755
rect 170 3710 220 3720
rect 480 3745 1380 3765
rect 480 3665 540 3745
rect 840 3665 890 3745
rect 910 3715 950 3725
rect 910 3695 920 3715
rect 940 3695 950 3715
rect 910 3685 950 3695
rect 480 3655 595 3665
rect 480 3635 490 3655
rect 530 3635 595 3655
rect 480 3625 595 3635
rect 840 3655 900 3665
rect 840 3635 850 3655
rect 890 3635 900 3655
rect 840 3625 900 3635
rect -175 3595 -125 3605
rect -175 3475 -165 3595
rect -135 3475 -125 3595
rect -175 3445 -125 3475
rect -55 3595 -5 3605
rect -55 3475 -45 3595
rect -15 3475 -5 3595
rect -55 3445 -5 3475
rect 65 3595 115 3605
rect 65 3475 75 3595
rect 105 3475 115 3595
rect 65 3445 115 3475
rect 185 3595 235 3605
rect 185 3475 195 3595
rect 225 3475 235 3595
rect 185 3445 235 3475
rect 305 3595 355 3605
rect 305 3475 315 3595
rect 345 3475 355 3595
rect 305 3465 355 3475
rect 425 3595 475 3605
rect 425 3475 435 3595
rect 465 3475 475 3595
rect -175 3435 300 3445
rect -175 3415 -165 3435
rect -70 3415 -45 3435
rect 50 3415 75 3435
rect 170 3415 195 3435
rect 290 3415 300 3435
rect -175 3405 300 3415
rect 425 3330 475 3475
rect 545 3595 595 3625
rect 920 3605 940 3685
rect 970 3665 1020 3745
rect 1320 3665 1380 3745
rect 1680 3745 1730 3755
rect 1680 3710 1690 3745
rect 1720 3710 1730 3745
rect 1680 3700 1730 3710
rect 960 3655 1020 3665
rect 960 3635 970 3655
rect 1010 3635 1020 3655
rect 960 3625 1020 3635
rect 1265 3655 1380 3665
rect 1265 3635 1330 3655
rect 1370 3635 1380 3655
rect 1265 3625 1380 3635
rect 545 3475 555 3595
rect 585 3475 595 3595
rect 545 3465 595 3475
rect 665 3595 715 3605
rect 665 3475 675 3595
rect 705 3475 715 3595
rect 665 3465 715 3475
rect 785 3595 835 3605
rect 785 3475 795 3595
rect 825 3475 835 3595
rect 785 3370 835 3475
rect 905 3595 955 3605
rect 905 3475 915 3595
rect 945 3475 955 3595
rect 905 3465 955 3475
rect 1025 3595 1075 3605
rect 1025 3475 1035 3595
rect 1065 3475 1075 3595
rect 1025 3370 1075 3475
rect 1145 3595 1195 3605
rect 1145 3475 1155 3595
rect 1185 3475 1195 3595
rect 1145 3465 1195 3475
rect 1265 3595 1315 3625
rect 1265 3475 1275 3595
rect 1305 3475 1315 3595
rect 1265 3465 1315 3475
rect 1385 3595 1435 3605
rect 1385 3475 1395 3595
rect 1425 3475 1435 3595
rect 785 3350 1075 3370
rect 1385 3330 1435 3475
rect 1505 3595 1555 3605
rect 1505 3475 1515 3595
rect 1545 3475 1555 3595
rect 1505 3465 1555 3475
rect 1625 3595 1675 3605
rect 1625 3475 1635 3595
rect 1665 3475 1675 3595
rect 1625 3445 1675 3475
rect 1745 3595 1795 3605
rect 1745 3475 1755 3595
rect 1785 3475 1795 3595
rect 1745 3445 1795 3475
rect 1865 3595 1915 3605
rect 1865 3475 1875 3595
rect 1905 3475 1915 3595
rect 1865 3445 1915 3475
rect 1985 3595 2035 3605
rect 1985 3475 1995 3595
rect 2025 3475 2035 3595
rect 1985 3445 2035 3475
rect 1560 3435 2035 3445
rect 1560 3415 1570 3435
rect 1665 3415 1690 3435
rect 1785 3415 1810 3435
rect 1905 3415 1930 3435
rect 2025 3415 2035 3435
rect 1560 3405 2035 3415
rect -225 3320 1435 3330
rect -225 3310 920 3320
rect 910 3300 920 3310
rect 940 3310 1435 3320
rect 940 3300 950 3310
rect 910 3290 950 3300
rect 2060 3290 2080 4175
rect 1030 3280 2080 3290
rect 1030 3260 1040 3280
rect 1060 3260 2080 3280
rect 1030 3250 2080 3260
rect 65 3210 1795 3230
rect -175 3100 -125 3110
rect -175 2980 -165 3100
rect -135 2980 -125 3100
rect -175 2950 -125 2980
rect -55 3100 -5 3110
rect -55 2980 -45 3100
rect -15 2980 -5 3100
rect -55 2970 -5 2980
rect 65 3100 115 3210
rect 65 2980 75 3100
rect 105 2980 115 3100
rect 65 2970 115 2980
rect 185 3100 235 3110
rect 185 2980 195 3100
rect 225 2980 235 3100
rect 185 2970 235 2980
rect 305 3100 355 3210
rect 305 2980 315 3100
rect 345 2980 355 3100
rect 305 2970 355 2980
rect 425 3180 475 3190
rect 425 3160 440 3180
rect 460 3160 475 3180
rect 425 3100 475 3160
rect 425 2980 435 3100
rect 465 2980 475 3100
rect -175 2940 -60 2950
rect -175 2920 -165 2940
rect -70 2920 -60 2940
rect -175 2910 -60 2920
rect 240 2870 350 2880
rect 240 2780 250 2870
rect 340 2780 350 2870
rect 425 2835 475 2980
rect 545 3100 595 3210
rect 545 2980 555 3100
rect 585 2980 595 3100
rect 545 2970 595 2980
rect 665 3100 715 3110
rect 665 2980 675 3100
rect 705 2980 715 3100
rect 665 2970 715 2980
rect 785 3100 835 3110
rect 785 2980 795 3100
rect 825 2980 835 3100
rect 785 2875 835 2980
rect 785 2850 795 2875
rect 825 2850 835 2875
rect 785 2840 835 2850
rect 905 3100 955 3110
rect 905 2980 915 3100
rect 945 2980 955 3100
rect 425 2810 435 2835
rect 465 2810 475 2835
rect 425 2800 475 2810
rect 240 2770 350 2780
rect 905 2755 955 2980
rect 1025 3100 1075 3110
rect 1025 2980 1035 3100
rect 1065 2980 1075 3100
rect 1025 2875 1075 2980
rect 1145 3100 1195 3110
rect 1145 2980 1155 3100
rect 1185 2980 1195 3100
rect 1145 2970 1195 2980
rect 1265 3100 1315 3210
rect 1265 2980 1275 3100
rect 1305 2980 1315 3100
rect 1265 2970 1315 2980
rect 1385 3100 1435 3110
rect 1385 2980 1395 3100
rect 1425 2980 1435 3100
rect 1025 2850 1035 2875
rect 1065 2850 1075 2875
rect 1025 2840 1075 2850
rect 1385 2835 1435 2980
rect 1505 3100 1555 3210
rect 1505 2980 1515 3100
rect 1545 2980 1555 3100
rect 1505 2970 1555 2980
rect 1625 3100 1675 3110
rect 1625 2980 1635 3100
rect 1665 2980 1675 3100
rect 1625 2970 1675 2980
rect 1745 3100 1795 3210
rect 1745 2980 1755 3100
rect 1785 2980 1795 3100
rect 1745 2970 1795 2980
rect 1865 3100 1915 3110
rect 1865 2980 1875 3100
rect 1905 2980 1915 3100
rect 1865 2970 1915 2980
rect 1985 3100 2035 3110
rect 1985 2980 1995 3100
rect 2025 2980 2035 3100
rect 1985 2950 2035 2980
rect 1920 2940 2035 2950
rect 1920 2920 1930 2940
rect 2025 2920 2035 2940
rect 1920 2910 2035 2920
rect 1385 2810 1395 2835
rect 1425 2810 1435 2835
rect 1385 2800 1435 2810
rect 1630 2870 1740 2880
rect 1630 2780 1640 2870
rect 1730 2780 1740 2870
rect 1630 2770 1740 2780
rect 460 2730 570 2740
rect 460 2640 470 2730
rect 560 2640 570 2730
rect 460 2630 570 2640
rect 665 2735 1195 2755
rect -175 2565 -125 2575
rect -175 2445 -165 2565
rect -135 2445 -125 2565
rect -175 2415 -125 2445
rect -55 2565 -5 2575
rect -55 2445 -45 2565
rect -15 2445 -5 2565
rect -55 2435 -5 2445
rect 65 2565 115 2575
rect 65 2445 75 2565
rect 105 2445 115 2565
rect -175 2405 -60 2415
rect -175 2385 -165 2405
rect -70 2385 -60 2405
rect -175 2375 -60 2385
rect 65 2335 115 2445
rect 185 2565 235 2575
rect 185 2445 195 2565
rect 225 2445 235 2565
rect 185 2435 235 2445
rect 305 2565 355 2575
rect 305 2445 315 2565
rect 345 2445 355 2565
rect 305 2335 355 2445
rect 425 2565 475 2575
rect 425 2445 435 2565
rect 465 2445 475 2565
rect 425 2435 475 2445
rect 545 2565 595 2575
rect 545 2445 555 2565
rect 585 2445 595 2565
rect 545 2335 595 2445
rect 665 2565 715 2735
rect 665 2445 675 2565
rect 705 2445 715 2565
rect 665 2435 715 2445
rect 785 2695 920 2705
rect 940 2695 1075 2705
rect 785 2685 1075 2695
rect 785 2565 835 2685
rect 785 2445 795 2565
rect 825 2445 835 2565
rect 785 2435 835 2445
rect 905 2655 955 2665
rect 905 2630 915 2655
rect 945 2630 955 2655
rect 905 2565 955 2630
rect 905 2445 915 2565
rect 945 2445 955 2565
rect 905 2435 955 2445
rect 1025 2565 1075 2685
rect 1025 2445 1035 2565
rect 1065 2445 1075 2565
rect 1025 2435 1075 2445
rect 1145 2565 1195 2735
rect 1305 2730 1415 2740
rect 1305 2640 1315 2730
rect 1405 2640 1415 2730
rect 1305 2630 1415 2640
rect 1145 2445 1155 2565
rect 1185 2445 1195 2565
rect 1145 2435 1195 2445
rect 1265 2565 1315 2575
rect 1265 2445 1275 2565
rect 1305 2445 1315 2565
rect 910 2385 950 2435
rect 910 2365 920 2385
rect 940 2365 950 2385
rect 910 2355 950 2365
rect 1265 2335 1315 2445
rect 1385 2565 1435 2575
rect 1385 2445 1395 2565
rect 1425 2445 1435 2565
rect 1385 2435 1435 2445
rect 1505 2565 1555 2575
rect 1505 2445 1515 2565
rect 1545 2445 1555 2565
rect 1505 2335 1555 2445
rect 1625 2565 1675 2575
rect 1625 2445 1635 2565
rect 1665 2445 1675 2565
rect 1625 2435 1675 2445
rect 1745 2565 1795 2575
rect 1745 2445 1755 2565
rect 1785 2445 1795 2565
rect 1745 2335 1795 2445
rect 1865 2565 1915 2575
rect 1865 2445 1875 2565
rect 1905 2445 1915 2565
rect 1865 2435 1915 2445
rect 1985 2565 2035 2575
rect 1985 2445 1995 2565
rect 2025 2445 2035 2565
rect 1985 2415 2035 2445
rect 1920 2405 2035 2415
rect 1920 2385 1930 2405
rect 2025 2385 2035 2405
rect 1920 2375 2035 2385
rect 65 2315 1795 2335
<< viali >>
rect 920 3300 940 3320
rect 1040 3260 1060 3280
rect 1035 2850 1065 2875
rect 920 2695 940 2715
<< metal1 >>
rect 910 3320 950 3330
rect 910 3300 920 3320
rect 940 3300 950 3320
rect 910 2715 950 3300
rect 1025 3280 1075 3295
rect 1025 3260 1040 3280
rect 1060 3260 1075 3280
rect 1025 2875 1075 3260
rect 1025 2850 1035 2875
rect 1065 2850 1075 2875
rect 1025 2840 1075 2850
rect 910 2695 920 2715
rect 940 2695 950 2715
rect 910 2685 950 2695
<< end >>
