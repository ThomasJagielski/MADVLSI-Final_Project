magic
tech sky130A
magscale 1 2
timestamp 1620714218
<< nwell >>
rect 4910 -4470 5590 -830
rect 4630 -5150 5590 -4470
rect 4910 -6210 5590 -5150
<< pwell >>
rect 3150 -187 3946 -34
rect 3150 -677 3303 -187
rect 3793 -677 3946 -187
rect 3150 -830 3946 -677
rect 3150 -1187 3946 -1034
rect 3150 -1677 3303 -1187
rect 3793 -1677 3946 -1187
rect 3150 -1830 3946 -1677
<< nbase >>
rect 3303 -677 3793 -187
rect 3303 -1677 3793 -1187
rect 2460 -3540 2540 -3440
<< pmos >>
rect 4950 -1230 5550 -1110
rect 4950 -1720 5550 -1600
rect 4950 -1960 5550 -1840
rect 4950 -2200 5550 -2080
rect 4950 -2440 5550 -2320
rect 4950 -2680 5550 -2560
rect 4950 -2920 5550 -2800
rect 4950 -3160 5550 -3040
rect 4950 -3400 5550 -3280
rect 4950 -3880 5550 -3760
rect 4950 -4120 5550 -4000
rect 4950 -4360 5550 -4240
rect 4950 -4600 5550 -4480
rect 4950 -4840 5550 -4720
rect 4950 -5080 5550 -4960
rect 4950 -5320 5550 -5200
rect 4950 -5560 5550 -5440
rect 4950 -6050 5550 -5930
<< pdiff >>
rect 3480 -381 3616 -364
rect 3480 -483 3497 -381
rect 3599 -483 3616 -381
rect 3480 -500 3616 -483
rect 4950 -1110 5550 -1000
rect 3480 -1381 3616 -1364
rect 3480 -1483 3497 -1381
rect 3599 -1483 3616 -1381
rect 3480 -1500 3616 -1483
rect 4950 -1370 5550 -1230
rect 4950 -1600 5550 -1480
rect 4950 -1840 5550 -1720
rect 4950 -2080 5550 -1960
rect 4950 -2320 5550 -2200
rect 4950 -2560 5550 -2440
rect 4950 -2800 5550 -2680
rect 4950 -3040 5550 -2920
rect 4950 -3280 5550 -3160
rect 4950 -3520 5550 -3400
rect 4950 -3760 5550 -3640
rect 4950 -4000 5550 -3880
rect 4950 -4240 5550 -4120
rect 4950 -4480 5550 -4360
rect 4950 -4720 5550 -4600
rect 4950 -4960 5550 -4840
rect 4950 -5200 5550 -5080
rect 4950 -5440 5550 -5320
rect 4950 -5690 5550 -5560
rect 4950 -5930 5550 -5800
rect 4950 -6170 5550 -6050
<< pdiffc >>
rect 3497 -483 3599 -381
rect 3497 -1483 3599 -1381
<< psubdiff >>
rect 3176 -94 3920 -60
rect 3176 -128 3210 -94
rect 3244 -128 3278 -94
rect 3312 -128 3346 -94
rect 3380 -128 3414 -94
rect 3448 -128 3648 -94
rect 3682 -128 3716 -94
rect 3750 -128 3784 -94
rect 3818 -128 3852 -94
rect 3886 -128 3920 -94
rect 3176 -161 3920 -128
rect 3176 -162 3277 -161
rect 3176 -196 3210 -162
rect 3244 -196 3277 -162
rect 3176 -230 3277 -196
rect 3819 -162 3920 -161
rect 3819 -196 3852 -162
rect 3886 -196 3920 -162
rect 3176 -264 3210 -230
rect 3244 -264 3277 -230
rect 3176 -298 3277 -264
rect 3176 -332 3210 -298
rect 3244 -332 3277 -298
rect 3176 -532 3277 -332
rect 3176 -566 3210 -532
rect 3244 -566 3277 -532
rect 3176 -600 3277 -566
rect 3176 -634 3210 -600
rect 3244 -634 3277 -600
rect 3176 -668 3277 -634
rect 3819 -230 3920 -196
rect 3819 -264 3852 -230
rect 3886 -264 3920 -230
rect 3819 -298 3920 -264
rect 3819 -332 3852 -298
rect 3886 -332 3920 -298
rect 3819 -532 3920 -332
rect 3819 -566 3852 -532
rect 3886 -566 3920 -532
rect 3819 -600 3920 -566
rect 3819 -634 3852 -600
rect 3886 -634 3920 -600
rect 3176 -702 3210 -668
rect 3244 -702 3277 -668
rect 3176 -703 3277 -702
rect 3819 -668 3920 -634
rect 3819 -702 3852 -668
rect 3886 -702 3920 -668
rect 3819 -703 3920 -702
rect 3176 -736 3920 -703
rect 3176 -770 3210 -736
rect 3244 -770 3278 -736
rect 3312 -770 3346 -736
rect 3380 -770 3414 -736
rect 3448 -770 3648 -736
rect 3682 -770 3716 -736
rect 3750 -770 3784 -736
rect 3818 -770 3852 -736
rect 3886 -770 3920 -736
rect 3176 -804 3920 -770
rect 3176 -1094 3920 -1060
rect 3176 -1128 3210 -1094
rect 3244 -1128 3278 -1094
rect 3312 -1128 3346 -1094
rect 3380 -1128 3414 -1094
rect 3448 -1128 3648 -1094
rect 3682 -1128 3716 -1094
rect 3750 -1128 3784 -1094
rect 3818 -1128 3852 -1094
rect 3886 -1128 3920 -1094
rect 3176 -1161 3920 -1128
rect 3176 -1162 3277 -1161
rect 3176 -1196 3210 -1162
rect 3244 -1196 3277 -1162
rect 3176 -1230 3277 -1196
rect 3819 -1162 3920 -1161
rect 3819 -1196 3852 -1162
rect 3886 -1196 3920 -1162
rect 3176 -1264 3210 -1230
rect 3244 -1264 3277 -1230
rect 3176 -1298 3277 -1264
rect 3176 -1332 3210 -1298
rect 3244 -1332 3277 -1298
rect 3176 -1532 3277 -1332
rect 3176 -1566 3210 -1532
rect 3244 -1566 3277 -1532
rect 3176 -1600 3277 -1566
rect 3176 -1634 3210 -1600
rect 3244 -1634 3277 -1600
rect 3176 -1668 3277 -1634
rect 3819 -1230 3920 -1196
rect 3819 -1264 3852 -1230
rect 3886 -1264 3920 -1230
rect 3819 -1298 3920 -1264
rect 3819 -1332 3852 -1298
rect 3886 -1332 3920 -1298
rect 3819 -1532 3920 -1332
rect 3819 -1566 3852 -1532
rect 3886 -1566 3920 -1532
rect 3819 -1600 3920 -1566
rect 3819 -1634 3852 -1600
rect 3886 -1634 3920 -1600
rect 3176 -1702 3210 -1668
rect 3244 -1702 3277 -1668
rect 3176 -1703 3277 -1702
rect 3819 -1668 3920 -1634
rect 3819 -1702 3852 -1668
rect 3886 -1702 3920 -1668
rect 3819 -1703 3920 -1702
rect 3176 -1736 3920 -1703
rect 3176 -1770 3210 -1736
rect 3244 -1770 3278 -1736
rect 3312 -1770 3346 -1736
rect 3380 -1770 3414 -1736
rect 3448 -1770 3648 -1736
rect 3682 -1770 3716 -1736
rect 3750 -1770 3784 -1736
rect 3818 -1770 3852 -1736
rect 3886 -1770 3920 -1736
rect 3176 -1804 3920 -1770
<< nsubdiff >>
rect 3339 -247 3757 -223
rect 3339 -281 3363 -247
rect 3397 -281 3431 -247
rect 3465 -281 3631 -247
rect 3665 -281 3699 -247
rect 3733 -281 3757 -247
rect 3339 -295 3757 -281
rect 3339 -315 3411 -295
rect 3339 -349 3363 -315
rect 3397 -349 3411 -315
rect 3339 -515 3411 -349
rect 3685 -315 3757 -295
rect 3685 -349 3699 -315
rect 3733 -349 3757 -315
rect 3339 -549 3363 -515
rect 3397 -549 3411 -515
rect 3339 -569 3411 -549
rect 3685 -515 3757 -349
rect 3685 -549 3699 -515
rect 3733 -549 3757 -515
rect 3685 -569 3757 -549
rect 3339 -583 3757 -569
rect 3339 -617 3363 -583
rect 3397 -617 3431 -583
rect 3465 -617 3631 -583
rect 3665 -617 3699 -583
rect 3733 -617 3757 -583
rect 3339 -641 3757 -617
rect 4950 -900 5550 -870
rect 4950 -980 4980 -900
rect 5520 -980 5550 -900
rect 4950 -1000 5550 -980
rect 3339 -1247 3757 -1223
rect 3339 -1281 3363 -1247
rect 3397 -1281 3431 -1247
rect 3465 -1281 3631 -1247
rect 3665 -1281 3699 -1247
rect 3733 -1281 3757 -1247
rect 3339 -1295 3757 -1281
rect 3339 -1315 3411 -1295
rect 3339 -1349 3363 -1315
rect 3397 -1349 3411 -1315
rect 3339 -1515 3411 -1349
rect 3685 -1315 3757 -1295
rect 3685 -1349 3699 -1315
rect 3733 -1349 3757 -1315
rect 3339 -1549 3363 -1515
rect 3397 -1549 3411 -1515
rect 3339 -1569 3411 -1549
rect 3685 -1515 3757 -1349
rect 3685 -1549 3699 -1515
rect 3733 -1549 3757 -1515
rect 3685 -1569 3757 -1549
rect 3339 -1583 3757 -1569
rect 3339 -1617 3363 -1583
rect 3397 -1617 3431 -1583
rect 3465 -1617 3631 -1583
rect 3665 -1617 3699 -1583
rect 3733 -1617 3757 -1583
rect 3339 -1641 3757 -1617
rect 4670 -4540 4800 -4510
rect 4670 -5080 4690 -4540
rect 4770 -5080 4800 -4540
rect 4670 -5110 4800 -5080
<< psubdiffcont >>
rect 3210 -128 3244 -94
rect 3278 -128 3312 -94
rect 3346 -128 3380 -94
rect 3414 -128 3448 -94
rect 3648 -128 3682 -94
rect 3716 -128 3750 -94
rect 3784 -128 3818 -94
rect 3852 -128 3886 -94
rect 3210 -196 3244 -162
rect 3852 -196 3886 -162
rect 3210 -264 3244 -230
rect 3210 -332 3244 -298
rect 3210 -566 3244 -532
rect 3210 -634 3244 -600
rect 3852 -264 3886 -230
rect 3852 -332 3886 -298
rect 3852 -566 3886 -532
rect 3852 -634 3886 -600
rect 3210 -702 3244 -668
rect 3852 -702 3886 -668
rect 3210 -770 3244 -736
rect 3278 -770 3312 -736
rect 3346 -770 3380 -736
rect 3414 -770 3448 -736
rect 3648 -770 3682 -736
rect 3716 -770 3750 -736
rect 3784 -770 3818 -736
rect 3852 -770 3886 -736
rect 3210 -1128 3244 -1094
rect 3278 -1128 3312 -1094
rect 3346 -1128 3380 -1094
rect 3414 -1128 3448 -1094
rect 3648 -1128 3682 -1094
rect 3716 -1128 3750 -1094
rect 3784 -1128 3818 -1094
rect 3852 -1128 3886 -1094
rect 3210 -1196 3244 -1162
rect 3852 -1196 3886 -1162
rect 3210 -1264 3244 -1230
rect 3210 -1332 3244 -1298
rect 3210 -1566 3244 -1532
rect 3210 -1634 3244 -1600
rect 3852 -1264 3886 -1230
rect 3852 -1332 3886 -1298
rect 3852 -1566 3886 -1532
rect 3852 -1634 3886 -1600
rect 3210 -1702 3244 -1668
rect 3852 -1702 3886 -1668
rect 3210 -1770 3244 -1736
rect 3278 -1770 3312 -1736
rect 3346 -1770 3380 -1736
rect 3414 -1770 3448 -1736
rect 3648 -1770 3682 -1736
rect 3716 -1770 3750 -1736
rect 3784 -1770 3818 -1736
rect 3852 -1770 3886 -1736
<< nsubdiffcont >>
rect 3363 -281 3397 -247
rect 3431 -281 3465 -247
rect 3631 -281 3665 -247
rect 3699 -281 3733 -247
rect 3363 -349 3397 -315
rect 3699 -349 3733 -315
rect 3363 -549 3397 -515
rect 3699 -549 3733 -515
rect 3363 -617 3397 -583
rect 3431 -617 3465 -583
rect 3631 -617 3665 -583
rect 3699 -617 3733 -583
rect 4980 -980 5520 -900
rect 3363 -1281 3397 -1247
rect 3431 -1281 3465 -1247
rect 3631 -1281 3665 -1247
rect 3699 -1281 3733 -1247
rect 3363 -1349 3397 -1315
rect 3699 -1349 3733 -1315
rect 3363 -1549 3397 -1515
rect 3699 -1549 3733 -1515
rect 3363 -1617 3397 -1583
rect 3431 -1617 3465 -1583
rect 3631 -1617 3665 -1583
rect 3699 -1617 3733 -1583
rect 4690 -5080 4770 -4540
<< poly >>
rect 15700 5820 15780 5840
rect 15700 5780 15720 5820
rect 15760 5790 15780 5820
rect 15760 5780 15820 5790
rect 15700 5760 15820 5780
rect -4290 5710 -4210 5730
rect -4290 5670 -4270 5710
rect -4230 5680 -4210 5710
rect 5730 5710 5810 5730
rect -4230 5670 -4170 5680
rect -4290 5650 -4170 5670
rect 5730 5670 5750 5710
rect 5790 5680 5810 5710
rect 5790 5670 5850 5680
rect 5730 5650 5850 5670
rect 15620 4320 15820 4340
rect 15620 4280 15640 4320
rect 15680 4310 15820 4320
rect 15680 4280 15700 4310
rect -4360 4260 -4280 4280
rect -4360 4220 -4340 4260
rect -4300 4230 -4280 4260
rect 5680 4260 5760 4280
rect 15620 4260 15700 4280
rect -4300 4220 -4140 4230
rect -4360 4200 -4140 4220
rect 5680 4220 5700 4260
rect 5740 4230 5760 4260
rect 5740 4220 5990 4230
rect 5680 4200 5990 4220
rect 5690 -1020 5980 -1000
rect 5690 -1060 5710 -1020
rect 5750 -1040 5980 -1020
rect 5750 -1060 5770 -1040
rect 5690 -1080 5770 -1060
rect 4890 -1230 4950 -1110
rect 5550 -1230 5580 -1110
rect 4890 -1600 4920 -1230
rect 4890 -1720 4950 -1600
rect 5550 -1720 5580 -1600
rect 4890 -1840 4920 -1720
rect 4890 -1960 4950 -1840
rect 5550 -1960 5580 -1840
rect 4890 -2080 4920 -1960
rect 4890 -2200 4950 -2080
rect 5550 -2200 5580 -2080
rect 4890 -2320 4920 -2200
rect 4890 -2440 4950 -2320
rect 5550 -2440 5580 -2320
rect 5770 -2430 5850 -2410
rect 4890 -2560 4920 -2440
rect 5770 -2470 5790 -2430
rect 5830 -2450 5850 -2430
rect 5830 -2470 5990 -2450
rect 5770 -2490 5990 -2470
rect 4890 -2680 4950 -2560
rect 5550 -2680 5580 -2560
rect 4890 -2800 4920 -2680
rect 4890 -2920 4950 -2800
rect 5550 -2920 5580 -2800
rect 4890 -3040 4920 -2920
rect 4890 -3160 4950 -3040
rect 5550 -3160 5580 -3040
rect 4890 -3280 4920 -3160
rect 4890 -3400 4950 -3280
rect 5550 -3400 5580 -3280
rect 4890 -3760 4920 -3400
rect 4890 -3880 4950 -3760
rect 5550 -3880 5580 -3760
rect 4890 -4000 4920 -3880
rect 4890 -4120 4950 -4000
rect 5550 -4120 5580 -4000
rect 4890 -4240 4920 -4120
rect 4890 -4360 4950 -4240
rect 5550 -4360 5580 -4240
rect 4890 -4480 4920 -4360
rect 4890 -4600 4950 -4480
rect 5550 -4600 5580 -4480
rect 4890 -4720 4920 -4600
rect 4890 -4840 4950 -4720
rect 5550 -4840 5580 -4720
rect 4890 -4960 4920 -4840
rect 4890 -5080 4950 -4960
rect 5550 -5080 5580 -4960
rect 4890 -5200 4920 -5080
rect 4890 -5320 4950 -5200
rect 5550 -5320 5580 -5200
rect 4890 -5440 4920 -5320
rect 4890 -5560 4950 -5440
rect 5550 -5560 5580 -5440
rect 4890 -5930 4920 -5560
rect 4860 -6050 4950 -5930
rect 5550 -6050 5580 -5930
rect 4860 -6240 4890 -6050
rect 4860 -6260 4940 -6240
rect 4860 -6300 4880 -6260
rect 4920 -6300 4940 -6260
rect 4860 -6320 4940 -6300
<< polycont >>
rect 15720 5780 15760 5820
rect -4270 5670 -4230 5710
rect 5750 5670 5790 5710
rect 15640 4280 15680 4320
rect -4340 4220 -4300 4260
rect 5700 4220 5740 4260
rect 5710 -1060 5750 -1020
rect 5790 -2470 5830 -2430
rect 4880 -6300 4920 -6260
<< locali >>
rect 15700 7160 21780 7200
rect -4290 6990 1790 7030
rect -4290 5730 -4250 6990
rect -4290 5710 -4210 5730
rect -4290 5670 -4270 5710
rect -4230 5670 -4210 5710
rect -4290 5650 -4210 5670
rect -4360 4260 -4280 4280
rect -4360 4220 -4340 4260
rect -4300 4220 -4280 4260
rect -4360 4200 -4280 4220
rect 1750 1590 1790 6990
rect 5730 6990 11800 7030
rect 5730 5730 5770 6990
rect 5730 5710 5810 5730
rect 5730 5670 5750 5710
rect 5790 5670 5810 5710
rect 5730 5650 5810 5670
rect 5680 4260 5760 4280
rect 5680 4220 5700 4260
rect 5740 4220 5760 4260
rect 5680 4200 5760 4220
rect 11760 1590 11800 6990
rect 15700 5840 15740 7160
rect 15700 5820 15780 5840
rect 15700 5780 15720 5820
rect 15760 5780 15780 5820
rect 15700 5760 15780 5780
rect 15620 4320 15700 4340
rect 15620 4280 15640 4320
rect 15680 4280 15700 4320
rect 15620 4260 15700 4280
rect 15620 200 15660 4260
rect 21740 1700 21780 7160
rect 4060 160 15660 200
rect 3176 -94 3920 -60
rect 3176 -128 3210 -94
rect 3244 -128 3278 -94
rect 3312 -128 3346 -94
rect 3380 -128 3414 -94
rect 3448 -128 3648 -94
rect 3682 -128 3716 -94
rect 3750 -128 3784 -94
rect 3818 -128 3852 -94
rect 3886 -128 3920 -94
rect 3176 -161 3920 -128
rect 3176 -162 3277 -161
rect 3176 -196 3210 -162
rect 3244 -196 3277 -162
rect 3176 -230 3277 -196
rect 3819 -162 3920 -161
rect 3819 -196 3852 -162
rect 3886 -196 3920 -162
rect 3176 -264 3210 -230
rect 3244 -264 3277 -230
rect 3176 -298 3277 -264
rect 3176 -332 3210 -298
rect 3244 -332 3277 -298
rect 3176 -532 3277 -332
rect 3176 -566 3210 -532
rect 3244 -566 3277 -532
rect 3176 -600 3277 -566
rect 3176 -634 3210 -600
rect 3244 -634 3277 -600
rect 3176 -668 3277 -634
rect 3339 -247 3757 -223
rect 3339 -281 3363 -247
rect 3397 -281 3431 -247
rect 3465 -281 3631 -247
rect 3665 -281 3699 -247
rect 3733 -281 3757 -247
rect 3339 -295 3757 -281
rect 3339 -315 3411 -295
rect 3339 -349 3363 -315
rect 3397 -349 3411 -315
rect 3339 -515 3411 -349
rect 3685 -315 3757 -295
rect 3685 -349 3699 -315
rect 3733 -349 3757 -315
rect 3469 -367 3627 -353
rect 3469 -401 3483 -367
rect 3517 -381 3579 -367
rect 3613 -401 3627 -367
rect 3469 -463 3497 -401
rect 3599 -463 3627 -401
rect 3469 -497 3483 -463
rect 3517 -497 3579 -483
rect 3613 -497 3627 -463
rect 3469 -511 3627 -497
rect 3339 -549 3363 -515
rect 3397 -549 3411 -515
rect 3339 -569 3411 -549
rect 3685 -515 3757 -349
rect 3685 -549 3699 -515
rect 3733 -549 3757 -515
rect 3685 -569 3757 -549
rect 3339 -583 3757 -569
rect 3339 -617 3363 -583
rect 3397 -617 3431 -583
rect 3465 -617 3631 -583
rect 3665 -617 3699 -583
rect 3733 -617 3757 -583
rect 3339 -641 3757 -617
rect 3819 -230 3920 -196
rect 3819 -264 3852 -230
rect 3886 -264 3920 -230
rect 3819 -298 3920 -264
rect 3819 -332 3852 -298
rect 3886 -332 3920 -298
rect 3819 -532 3920 -332
rect 3819 -566 3852 -532
rect 3886 -566 3920 -532
rect 3819 -600 3920 -566
rect 3819 -634 3852 -600
rect 3886 -634 3920 -600
rect 3176 -702 3210 -668
rect 3244 -702 3277 -668
rect 3176 -703 3277 -702
rect 3819 -668 3920 -634
rect 3819 -702 3852 -668
rect 3886 -702 3920 -668
rect 3819 -703 3920 -702
rect 3176 -736 3920 -703
rect 3176 -770 3210 -736
rect 3244 -770 3278 -736
rect 3312 -770 3346 -736
rect 3380 -770 3414 -736
rect 3448 -770 3648 -736
rect 3682 -770 3716 -736
rect 3750 -770 3784 -736
rect 3818 -770 3852 -736
rect 3886 -770 3920 -736
rect 3176 -804 3920 -770
rect 1820 -1160 2360 -1060
rect 3176 -1094 3920 -1060
rect 3176 -1128 3210 -1094
rect 3244 -1128 3278 -1094
rect 3312 -1128 3346 -1094
rect 3380 -1128 3414 -1094
rect 3448 -1128 3648 -1094
rect 3682 -1128 3716 -1094
rect 3750 -1128 3784 -1094
rect 3818 -1128 3852 -1094
rect 3886 -1128 3920 -1094
rect 3176 -1161 3920 -1128
rect 3176 -1162 3277 -1161
rect 3176 -1196 3210 -1162
rect 3244 -1196 3277 -1162
rect 1690 -1300 2410 -1220
rect 3176 -1230 3277 -1196
rect 3819 -1162 3920 -1161
rect 3819 -1196 3852 -1162
rect 3886 -1196 3920 -1162
rect 3176 -1264 3210 -1230
rect 3244 -1264 3277 -1230
rect 3176 -1298 3277 -1264
rect 3176 -1332 3210 -1298
rect 3244 -1332 3277 -1298
rect 3176 -1532 3277 -1332
rect 3176 -1566 3210 -1532
rect 3244 -1566 3277 -1532
rect 3176 -1600 3277 -1566
rect 3176 -1634 3210 -1600
rect 3244 -1634 3277 -1600
rect 3176 -1668 3277 -1634
rect 3339 -1247 3757 -1223
rect 3339 -1281 3363 -1247
rect 3397 -1281 3431 -1247
rect 3465 -1281 3631 -1247
rect 3665 -1281 3699 -1247
rect 3733 -1281 3757 -1247
rect 3339 -1295 3757 -1281
rect 3339 -1315 3411 -1295
rect 3339 -1349 3363 -1315
rect 3397 -1349 3411 -1315
rect 3339 -1515 3411 -1349
rect 3685 -1315 3757 -1295
rect 3685 -1349 3699 -1315
rect 3733 -1349 3757 -1315
rect 3469 -1367 3627 -1353
rect 3469 -1401 3483 -1367
rect 3517 -1381 3579 -1367
rect 3613 -1401 3627 -1367
rect 3469 -1463 3497 -1401
rect 3599 -1463 3627 -1401
rect 3469 -1497 3483 -1463
rect 3517 -1497 3579 -1483
rect 3613 -1497 3627 -1463
rect 3469 -1511 3627 -1497
rect 3339 -1549 3363 -1515
rect 3397 -1549 3411 -1515
rect 3339 -1569 3411 -1549
rect 3685 -1515 3757 -1349
rect 3685 -1549 3699 -1515
rect 3733 -1549 3757 -1515
rect 3685 -1569 3757 -1549
rect 3339 -1583 3757 -1569
rect 3339 -1617 3363 -1583
rect 3397 -1617 3431 -1583
rect 3465 -1617 3631 -1583
rect 3665 -1617 3699 -1583
rect 3733 -1617 3757 -1583
rect 3339 -1641 3757 -1617
rect 3819 -1230 3920 -1196
rect 3819 -1264 3852 -1230
rect 3886 -1264 3920 -1230
rect 3819 -1298 3920 -1264
rect 3819 -1332 3852 -1298
rect 3886 -1332 3920 -1298
rect 3819 -1532 3920 -1332
rect 3819 -1566 3852 -1532
rect 3886 -1566 3920 -1532
rect 3819 -1600 3920 -1566
rect 3819 -1634 3852 -1600
rect 3886 -1634 3920 -1600
rect 3176 -1702 3210 -1668
rect 3244 -1702 3277 -1668
rect 3176 -1703 3277 -1702
rect 3819 -1668 3920 -1634
rect 3819 -1702 3852 -1668
rect 3886 -1702 3920 -1668
rect 3819 -1703 3920 -1702
rect 3176 -1736 3920 -1703
rect 3176 -1770 3210 -1736
rect 3244 -1770 3278 -1736
rect 3312 -1770 3346 -1736
rect 3380 -1770 3414 -1736
rect 3448 -1770 3648 -1736
rect 3682 -1770 3716 -1736
rect 3750 -1770 3784 -1736
rect 3818 -1770 3852 -1736
rect 3886 -1770 3920 -1736
rect 3176 -1804 3920 -1770
rect 4060 -1950 4100 160
rect 4960 -900 5540 -880
rect 4960 -980 4980 -900
rect 5520 -980 5540 -900
rect 4960 -1020 5540 -980
rect 4960 -1080 4980 -1020
rect 5520 -1080 5540 -1020
rect 4960 -1100 5540 -1080
rect 5690 -1020 5770 -1000
rect 5690 -1060 5710 -1020
rect 5750 -1060 5770 -1020
rect 5690 -1080 5770 -1060
rect 4960 -1260 5540 -1250
rect 4960 -1340 4980 -1260
rect 5520 -1340 5540 -1260
rect 4960 -1350 5540 -1340
rect 4870 -1590 5540 -1480
rect 4870 -1950 4910 -1590
rect 4960 -1830 5630 -1730
rect 2610 -1970 4910 -1950
rect 2610 -1990 5540 -1970
rect 2810 -2160 2920 -2060
rect 4870 -2070 5540 -1990
rect 4870 -2450 4910 -2070
rect 5590 -2210 5630 -1830
rect 4960 -2310 5630 -2210
rect 4870 -2550 5540 -2450
rect 4870 -2930 4910 -2550
rect 5590 -2690 5630 -2310
rect 4960 -2790 5630 -2690
rect 4870 -3030 5540 -2930
rect 4870 -3410 4910 -3030
rect 5590 -3170 5630 -2790
rect 4960 -3270 5630 -3170
rect 5690 -3310 5730 -1080
rect 5590 -3350 5730 -3310
rect 5770 -2430 5850 -2410
rect 5770 -2470 5790 -2430
rect 5830 -2470 5850 -2430
rect 5770 -2490 5850 -2470
rect 4870 -3510 5540 -3410
rect 4870 -3750 5540 -3650
rect 4870 -4130 4910 -3750
rect 5590 -3890 5630 -3350
rect 4960 -3990 5630 -3890
rect 4870 -4230 5540 -4130
rect 4670 -4540 4790 -4520
rect 2020 -5090 3930 -5050
rect 2020 -5200 2460 -5090
rect 3890 -6060 3930 -5090
rect 4670 -5080 4690 -4540
rect 4770 -5080 4790 -4540
rect 4670 -5100 4790 -5080
rect 4870 -4610 4910 -4230
rect 5590 -4370 5630 -3990
rect 4960 -4390 5630 -4370
rect 4960 -4450 4980 -4390
rect 5520 -4450 5630 -4390
rect 4960 -4470 5630 -4450
rect 4870 -4710 5540 -4610
rect 4870 -5090 4910 -4710
rect 5590 -4850 5630 -4470
rect 4960 -4950 5630 -4850
rect 4870 -5190 5540 -5090
rect 4870 -5570 4910 -5190
rect 5590 -5330 5630 -4950
rect 4960 -5430 5630 -5330
rect 4870 -5590 5540 -5570
rect 4870 -5660 4970 -5590
rect 5510 -5660 5540 -5590
rect 4870 -5670 5540 -5660
rect 4960 -5680 5540 -5670
rect 4960 -5830 5540 -5810
rect 4960 -5900 4980 -5830
rect 5520 -5900 5540 -5830
rect 4960 -5920 5540 -5900
rect 5770 -6060 5820 -2490
rect 3890 -6160 5820 -6060
rect 4860 -6260 4940 -6240
rect 4860 -6300 4880 -6260
rect 4920 -6280 4940 -6260
rect 11840 -6280 11880 -5050
rect 4920 -6300 11880 -6280
rect 4860 -6320 11880 -6300
<< viali >>
rect -4340 4220 -4300 4260
rect 5700 4220 5740 4260
rect 3483 -381 3517 -367
rect 3579 -381 3613 -367
rect 3483 -401 3497 -381
rect 3497 -401 3517 -381
rect 3579 -401 3599 -381
rect 3599 -401 3613 -381
rect 3483 -483 3497 -463
rect 3497 -483 3517 -463
rect 3579 -483 3599 -463
rect 3599 -483 3613 -463
rect 3483 -497 3517 -483
rect 3579 -497 3613 -483
rect 3483 -1381 3517 -1367
rect 3579 -1381 3613 -1367
rect 3483 -1401 3497 -1381
rect 3497 -1401 3517 -1381
rect 3579 -1401 3599 -1381
rect 3599 -1401 3613 -1381
rect 3483 -1483 3497 -1463
rect 3497 -1483 3517 -1463
rect 3579 -1483 3599 -1463
rect 3599 -1483 3613 -1463
rect 3483 -1497 3517 -1483
rect 3579 -1497 3613 -1483
rect 4980 -980 5520 -900
rect 4980 -1080 5520 -1020
rect 4980 -1340 5520 -1260
rect 2570 -1990 2610 -1950
rect 4690 -5080 4770 -4540
rect 4980 -4450 5520 -4390
rect 4970 -5660 5510 -5590
rect 4980 -5900 5520 -5830
<< metal1 >>
rect -4360 4260 -4280 4280
rect -4360 4220 -4340 4260
rect -4300 4220 -4280 4260
rect -4360 4200 -4280 4220
rect 5680 4260 5760 4280
rect 5680 4220 5700 4260
rect 5740 4220 5760 4260
rect 5680 4200 5760 4220
rect -4320 370 -4280 4200
rect 5720 370 5760 4200
rect -4320 330 5760 370
rect 3465 -367 3631 -349
rect 3465 -401 3483 -367
rect 3517 -401 3579 -367
rect 3613 -401 3631 -367
rect 3465 -463 3631 -401
rect 3465 -497 3483 -463
rect 3517 -497 3579 -463
rect 3613 -497 3631 -463
rect 3465 -515 3631 -497
rect 4000 -860 4160 330
rect 1470 -1020 4160 -860
rect 1470 -1350 1620 -1020
rect 4000 -1250 4160 -1020
rect 4950 -900 5550 -870
rect 4950 -980 4980 -900
rect 5520 -980 5550 -900
rect 4950 -990 5550 -980
rect 4950 -1020 5660 -990
rect 4950 -1080 4980 -1020
rect 5520 -1080 5660 -1020
rect 4950 -1110 5660 -1080
rect 4000 -1260 5540 -1250
rect 4000 -1340 4980 -1260
rect 5520 -1340 5540 -1260
rect 1470 -1490 2630 -1350
rect 1490 -1510 2630 -1490
rect 3465 -1367 3631 -1349
rect 4000 -1350 5540 -1340
rect 3465 -1401 3483 -1367
rect 3517 -1401 3579 -1367
rect 3613 -1401 3631 -1367
rect 3465 -1463 3631 -1401
rect 3465 -1497 3483 -1463
rect 3517 -1497 3579 -1463
rect 3613 -1497 3631 -1463
rect 3465 -1515 3631 -1497
rect 2550 -1950 2630 -1930
rect 2550 -1990 2570 -1950
rect 2610 -1990 2630 -1950
rect 2550 -2430 2630 -1990
rect 2460 -3450 2540 -3440
rect 2460 -3510 2470 -3450
rect 2530 -3510 2540 -3450
rect 2460 -3520 2540 -3510
rect 5880 -3680 6020 -3330
rect 4190 -3820 6020 -3680
rect 4960 -4390 5550 -4370
rect 4960 -4450 4980 -4390
rect 5520 -4450 5550 -4390
rect 4960 -4470 5550 -4450
rect 4670 -4540 4800 -4510
rect 4670 -5080 4690 -4540
rect 4770 -5080 4800 -4540
rect 4670 -5110 4800 -5080
rect 3719 -5210 5782 -5208
rect 3719 -5310 6720 -5210
rect 3719 -5311 5782 -5310
rect 3720 -5380 3820 -5311
rect 2970 -5480 3820 -5380
rect 4960 -5590 5540 -5570
rect 4960 -5660 4970 -5590
rect 5510 -5660 5540 -5590
rect 4960 -5680 5540 -5660
rect 4960 -5830 5540 -5810
rect 4960 -5900 4980 -5830
rect 5520 -5900 5540 -5830
rect 4960 -5920 5540 -5900
<< via1 >>
rect 4980 -980 5520 -900
rect 4980 -1080 5520 -1020
rect 2470 -3510 2530 -3450
rect 4980 -4450 5520 -4390
rect 4690 -5080 4770 -4540
rect 4970 -5660 5510 -5590
rect 4980 -5900 5520 -5830
<< metal2 >>
rect 4950 -900 5550 -870
rect 4950 -980 4980 -900
rect 5520 -980 5550 -900
rect 4950 -990 5550 -980
rect 4950 -1020 5660 -990
rect 4950 -1080 4980 -1020
rect 5520 -1080 5660 -1020
rect 4950 -1110 5660 -1080
rect 5620 -1230 5660 -1110
rect 5620 -1290 6140 -1230
rect 2460 -3450 2540 -3440
rect 2460 -3510 2470 -3450
rect 2530 -3510 2540 -3450
rect 2460 -3980 2540 -3510
rect 2460 -4020 4190 -3980
rect 4150 -4350 4190 -4020
rect 4150 -4390 5550 -4350
rect 4960 -4450 4980 -4390
rect 5520 -4450 5550 -4390
rect 4960 -4470 5550 -4450
rect 4670 -4540 4800 -4510
rect 4670 -5080 4690 -4540
rect 4770 -5080 4800 -4540
rect 4670 -5110 4800 -5080
rect 4960 -5590 5540 -5570
rect 4960 -5660 4970 -5590
rect 5510 -5660 5540 -5590
rect 4960 -5810 5540 -5660
rect 4960 -5830 5670 -5810
rect 4960 -5900 4980 -5830
rect 5520 -5900 5670 -5830
rect 4960 -5910 5670 -5900
rect 4960 -5920 5540 -5910
rect 5610 -6210 5670 -5910
rect 6370 -6210 6470 -5720
rect 5610 -6260 6470 -6210
<< comment >>
rect 3176 -47 3177 -34
tri 3177 -47 3181 -43 se
tri 3915 -47 3919 -43 sw
rect 3919 -47 3920 -34
rect 3176 -48 3521 -47
rect 3574 -48 3920 -47
rect 3176 -60 3177 -48
tri 3177 -52 3181 -48 ne
tri 3915 -52 3919 -48 nw
rect 3919 -60 3920 -48
rect 3303 -210 3304 -197
tri 3304 -210 3308 -206 se
tri 3788 -210 3792 -206 sw
rect 3792 -210 3793 -197
rect 3303 -211 3495 -210
rect 3602 -211 3793 -210
rect 3303 -223 3304 -211
tri 3304 -215 3308 -211 ne
tri 3788 -215 3792 -211 nw
rect 3792 -223 3793 -211
rect 3339 -265 3340 -252
tri 3340 -265 3344 -261 se
tri 3358 -265 3362 -261 sw
rect 3362 -265 3363 -252
rect 3339 -266 3363 -265
rect 3339 -278 3340 -266
tri 3340 -270 3344 -266 ne
tri 3349 -270 3351 -267 se
tri 3358 -270 3362 -266 nw
tri 3348 -273 3349 -270 se
rect 3349 -273 3351 -270
tri 3351 -273 3352 -270 sw
rect 3347 -274 3348 -273
tri 3348 -274 3349 -273 nw
rect 3351 -274 3352 -273
rect 3345 -306 3350 -274
rect 3362 -278 3363 -266
rect 3757 -297 3758 -284
tri 3758 -297 3762 -293 se
tri 3814 -297 3818 -293 sw
rect 3818 -297 3819 -284
rect 3757 -298 3819 -297
rect 3757 -310 3758 -298
tri 3758 -302 3762 -298 ne
tri 3814 -302 3818 -298 nw
rect 3818 -310 3819 -298
rect 3480 -351 3481 -338
tri 3481 -351 3485 -347 se
tri 3611 -351 3615 -347 sw
rect 3615 -351 3616 -338
rect 3480 -352 3527 -351
rect 3569 -352 3616 -351
rect 3480 -364 3481 -352
tri 3481 -356 3485 -352 ne
tri 3611 -356 3615 -352 nw
rect 3615 -364 3616 -352
rect 3339 -388 3340 -375
tri 3340 -388 3344 -384 se
tri 3406 -388 3410 -384 sw
rect 3410 -388 3411 -375
rect 3339 -389 3411 -388
rect 3339 -401 3340 -389
tri 3340 -393 3344 -389 ne
tri 3406 -393 3410 -389 nw
rect 3410 -401 3411 -389
tri 3540 -426 3542 -424 se
tri 3542 -426 3543 -424 sw
tri 3553 -426 3554 -424 se
tri 3554 -426 3556 -424 sw
tri 3540 -427 3542 -426 ne
rect 3542 -427 3543 -426
tri 3543 -427 3545 -426 sw
tri 3551 -427 3553 -426 se
tri 3542 -430 3545 -427 ne
tri 3545 -429 3546 -427 sw
tri 3550 -429 3551 -427 se
rect 3551 -429 3553 -427
tri 3553 -429 3556 -426 nw
rect 3545 -430 3546 -429
tri 3546 -430 3548 -429 sw
tri 3548 -430 3550 -429 se
tri 3545 -432 3546 -430 ne
tri 3543 -435 3546 -432 se
rect 3546 -434 3550 -430
tri 3550 -432 3553 -429 nw
rect 3546 -435 3547 -434
tri 3547 -435 3548 -434 nw
tri 3548 -435 3549 -434 ne
rect 3549 -435 3550 -434
tri 3550 -435 3553 -432 sw
tri 3540 -438 3543 -435 se
tri 3543 -438 3546 -435 nw
tri 3550 -438 3553 -435 ne
tri 3553 -438 3556 -435 sw
tri 3540 -440 3542 -438 ne
tri 3542 -440 3543 -438 nw
tri 3553 -440 3554 -438 ne
tri 3554 -440 3556 -438 nw
rect 3616 -500 3617 -487
tri 3617 -500 3621 -496 se
tri 3680 -500 3684 -496 sw
rect 3684 -500 3685 -487
rect 3616 -501 3685 -500
rect 3616 -513 3617 -501
tri 3617 -505 3621 -501 ne
tri 3680 -505 3684 -501 nw
rect 3684 -513 3685 -501
rect 3819 -500 3820 -487
tri 3820 -500 3824 -496 se
tri 3915 -500 3919 -496 sw
rect 3919 -500 3920 -487
rect 3819 -501 3920 -500
rect 3819 -513 3820 -501
tri 3820 -505 3824 -501 ne
tri 3915 -505 3919 -501 nw
rect 3919 -513 3920 -501
rect 3339 -654 3340 -641
tri 3340 -654 3344 -650 se
tri 3752 -654 3756 -650 sw
rect 3756 -654 3757 -641
rect 3339 -655 3527 -654
rect 3569 -655 3757 -654
rect 3339 -667 3340 -655
tri 3340 -659 3344 -655 ne
tri 3752 -659 3756 -655 nw
rect 3756 -667 3757 -655
rect 3512 -694 3513 -681
tri 3513 -694 3517 -690 se
tri 3579 -694 3583 -690 sw
rect 3583 -694 3584 -681
rect 3512 -695 3584 -694
rect 3512 -707 3513 -695
tri 3513 -699 3517 -695 ne
tri 3579 -699 3583 -695 nw
rect 3583 -707 3584 -695
rect 3176 -1047 3177 -1034
tri 3177 -1047 3181 -1043 se
tri 3915 -1047 3919 -1043 sw
rect 3919 -1047 3920 -1034
rect 3176 -1048 3521 -1047
rect 3574 -1048 3920 -1047
rect 3176 -1060 3177 -1048
tri 3177 -1052 3181 -1048 ne
tri 3915 -1052 3919 -1048 nw
rect 3919 -1060 3920 -1048
rect 3303 -1210 3304 -1197
tri 3304 -1210 3308 -1206 se
tri 3788 -1210 3792 -1206 sw
rect 3792 -1210 3793 -1197
rect 3303 -1211 3495 -1210
rect 3602 -1211 3793 -1210
rect 3303 -1223 3304 -1211
tri 3304 -1215 3308 -1211 ne
tri 3788 -1215 3792 -1211 nw
rect 3792 -1223 3793 -1211
rect 3339 -1265 3340 -1252
tri 3340 -1265 3344 -1261 se
tri 3358 -1265 3362 -1261 sw
rect 3362 -1265 3363 -1252
rect 3339 -1266 3363 -1265
rect 3339 -1278 3340 -1266
tri 3340 -1270 3344 -1266 ne
tri 3349 -1270 3351 -1267 se
tri 3358 -1270 3362 -1266 nw
tri 3348 -1273 3349 -1270 se
rect 3349 -1273 3351 -1270
tri 3351 -1273 3352 -1270 sw
rect 3347 -1274 3348 -1273
tri 3348 -1274 3349 -1273 nw
rect 3351 -1274 3352 -1273
rect 3345 -1306 3350 -1274
rect 3362 -1278 3363 -1266
rect 3757 -1297 3758 -1284
tri 3758 -1297 3762 -1293 se
tri 3814 -1297 3818 -1293 sw
rect 3818 -1297 3819 -1284
rect 3757 -1298 3819 -1297
rect 3757 -1310 3758 -1298
tri 3758 -1302 3762 -1298 ne
tri 3814 -1302 3818 -1298 nw
rect 3818 -1310 3819 -1298
rect 3480 -1351 3481 -1338
tri 3481 -1351 3485 -1347 se
tri 3611 -1351 3615 -1347 sw
rect 3615 -1351 3616 -1338
rect 3480 -1352 3527 -1351
rect 3569 -1352 3616 -1351
rect 3480 -1364 3481 -1352
tri 3481 -1356 3485 -1352 ne
tri 3611 -1356 3615 -1352 nw
rect 3615 -1364 3616 -1352
rect 3339 -1388 3340 -1375
tri 3340 -1388 3344 -1384 se
tri 3406 -1388 3410 -1384 sw
rect 3410 -1388 3411 -1375
rect 3339 -1389 3411 -1388
rect 3339 -1401 3340 -1389
tri 3340 -1393 3344 -1389 ne
tri 3406 -1393 3410 -1389 nw
rect 3410 -1401 3411 -1389
tri 3540 -1426 3542 -1424 se
tri 3542 -1426 3543 -1424 sw
tri 3553 -1426 3554 -1424 se
tri 3554 -1426 3556 -1424 sw
tri 3540 -1427 3542 -1426 ne
rect 3542 -1427 3543 -1426
tri 3543 -1427 3545 -1426 sw
tri 3551 -1427 3553 -1426 se
tri 3542 -1430 3545 -1427 ne
tri 3545 -1429 3546 -1427 sw
tri 3550 -1429 3551 -1427 se
rect 3551 -1429 3553 -1427
tri 3553 -1429 3556 -1426 nw
rect 3545 -1430 3546 -1429
tri 3546 -1430 3548 -1429 sw
tri 3548 -1430 3550 -1429 se
tri 3545 -1432 3546 -1430 ne
tri 3543 -1435 3546 -1432 se
rect 3546 -1434 3550 -1430
tri 3550 -1432 3553 -1429 nw
rect 3546 -1435 3547 -1434
tri 3547 -1435 3548 -1434 nw
tri 3548 -1435 3549 -1434 ne
rect 3549 -1435 3550 -1434
tri 3550 -1435 3553 -1432 sw
tri 3540 -1438 3543 -1435 se
tri 3543 -1438 3546 -1435 nw
tri 3550 -1438 3553 -1435 ne
tri 3553 -1438 3556 -1435 sw
tri 3540 -1440 3542 -1438 ne
tri 3542 -1440 3543 -1438 nw
tri 3553 -1440 3554 -1438 ne
tri 3554 -1440 3556 -1438 nw
rect 3616 -1500 3617 -1487
tri 3617 -1500 3621 -1496 se
tri 3680 -1500 3684 -1496 sw
rect 3684 -1500 3685 -1487
rect 3616 -1501 3685 -1500
rect 3616 -1513 3617 -1501
tri 3617 -1505 3621 -1501 ne
tri 3680 -1505 3684 -1501 nw
rect 3684 -1513 3685 -1501
rect 3819 -1500 3820 -1487
tri 3820 -1500 3824 -1496 se
tri 3915 -1500 3919 -1496 sw
rect 3919 -1500 3920 -1487
rect 3819 -1501 3920 -1500
rect 3819 -1513 3820 -1501
tri 3820 -1505 3824 -1501 ne
tri 3915 -1505 3919 -1501 nw
rect 3919 -1513 3920 -1501
rect 3339 -1654 3340 -1641
tri 3340 -1654 3344 -1650 se
tri 3752 -1654 3756 -1650 sw
rect 3756 -1654 3757 -1641
rect 3339 -1655 3527 -1654
rect 3569 -1655 3757 -1654
rect 3339 -1667 3340 -1655
tri 3340 -1659 3344 -1655 ne
tri 3752 -1659 3756 -1655 nw
rect 3756 -1667 3757 -1655
rect 3512 -1694 3513 -1681
tri 3513 -1694 3517 -1690 se
tri 3579 -1694 3583 -1690 sw
rect 3583 -1694 3584 -1681
rect 3512 -1695 3584 -1694
rect 3512 -1707 3513 -1695
tri 3513 -1699 3517 -1695 ne
tri 3579 -1699 3583 -1695 nw
rect 3583 -1707 3584 -1695
use bandgap_pnp  bandgap_pnp_0
timestamp 1620714017
transform 1 0 2150 0 1 -1830
box -4000 -4480 2310 1796
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620692581
transform 1 0 6478 0 1 -10866
box -510 4630 8890 10940
use selfbiasedcascode2stage  selfbiasedcascode2stage_1
timestamp 1620692581
transform 1 0 6340 0 1 -4180
box -510 4630 8890 10940
use selfbiasedcascode2stage  selfbiasedcascode2stage_2
timestamp 1620692581
transform 1 0 -3670 0 1 -4180
box -510 4630 8890 10940
use selfbiasedcascode2stage  selfbiasedcascode2stage_3
timestamp 1620692581
transform 1 0 16320 0 1 -4070
box -510 4630 8890 10940
<< labels >>
flabel locali s 3525 -452 3571 -408 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 3852 -447 3893 -421 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 3706 -446 3733 -420 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 3555 -740 3555 -740 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 3555 -607 3555 -607 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 3319 -313 3319 -313 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 3319 -334 3319 -334 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 3547 -682 3547 -682 0 FreeSans 100 0 0 0 0.360
flabel comment s 3548 -46 3548 -46 0 FreeSans 100 0 0 0 3.720
flabel comment s 3548 -209 3548 -209 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 3869 -488 3869 -488 0 FreeSans 100 0 0 0 0.505
flabel comment s 3788 -285 3788 -285 0 FreeSans 100 0 0 0 0.310
flabel comment s 3374 -376 3374 -376 0 FreeSans 100 0 0 0 0.360
flabel comment s 3650 -488 3650 -488 0 FreeSans 100 0 0 0 0.345
flabel comment s 3548 -653 3548 -653 0 FreeSans 100 0 0 0 2.090
flabel comment s 3548 -350 3548 -350 0 FreeSans 100 0 0 0 0.068
flabel locali s 3525 -1452 3571 -1408 0 FreeSans 200 0 0 0 Emitter
port 3 nsew
flabel locali s 3852 -1447 3893 -1421 0 FreeSans 200 0 0 0 Collector
port 2 nsew
flabel locali s 3706 -1446 3733 -1420 0 FreeSans 200 0 0 0 Base
port 1 nsew
flabel comment s 3555 -1740 3555 -1740 0 FreeSans 180 0 0 0 Use 28 licons in collector to match PNP model
flabel comment s 3555 -1607 3555 -1607 0 FreeSans 140 0 0 0 Use 12 licons in base to match PNP model
flabel comment s 3319 -1313 3319 -1313 0 FreeSans 100 0 0 0 0.12 min
flabel comment s 3319 -1334 3319 -1334 0 FreeSans 100 0 0 0 adj. sides
flabel comment s 3547 -1682 3547 -1682 0 FreeSans 100 0 0 0 0.360
flabel comment s 3548 -1046 3548 -1046 0 FreeSans 100 0 0 0 3.720
flabel comment s 3548 -1209 3548 -1209 0 FreeSans 100 0 0 0 2.450(nwell)
flabel comment s 3869 -1488 3869 -1488 0 FreeSans 100 0 0 0 0.505
flabel comment s 3788 -1285 3788 -1285 0 FreeSans 100 0 0 0 0.310
flabel comment s 3374 -1376 3374 -1376 0 FreeSans 100 0 0 0 0.360
flabel comment s 3650 -1488 3650 -1488 0 FreeSans 100 0 0 0 0.345
flabel comment s 3548 -1653 3548 -1653 0 FreeSans 100 0 0 0 2.090
flabel comment s 3548 -1350 3548 -1350 0 FreeSans 100 0 0 0 0.068
<< end >>
