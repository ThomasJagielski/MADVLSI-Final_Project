magic
tech sky130A
magscale 1 2
timestamp 1620719426
<< nwell >>
rect 4910 -4470 5590 -830
rect 4630 -5150 5590 -4470
rect 4910 -6210 5590 -5150
<< pmos >>
rect 4950 -1230 5550 -1110
rect 4950 -1720 5550 -1600
rect 4950 -1960 5550 -1840
rect 4950 -2200 5550 -2080
rect 4950 -2440 5550 -2320
rect 4950 -2680 5550 -2560
rect 4950 -2920 5550 -2800
rect 4950 -3160 5550 -3040
rect 4950 -3400 5550 -3280
rect 4950 -3880 5550 -3760
rect 4950 -4120 5550 -4000
rect 4950 -4360 5550 -4240
rect 4950 -4600 5550 -4480
rect 4950 -4840 5550 -4720
rect 4950 -5080 5550 -4960
rect 4950 -5320 5550 -5200
rect 4950 -5560 5550 -5440
rect 4950 -6050 5550 -5930
<< pdiff >>
rect 4950 -1110 5550 -1000
rect 4950 -1370 5550 -1230
rect 4950 -1600 5550 -1480
rect 4950 -1840 5550 -1720
rect 4950 -2080 5550 -1960
rect 4950 -2320 5550 -2200
rect 4950 -2560 5550 -2440
rect 4950 -2800 5550 -2680
rect 4950 -3040 5550 -2920
rect 4950 -3280 5550 -3160
rect 4950 -3520 5550 -3400
rect 4950 -3760 5550 -3640
rect 4950 -4000 5550 -3880
rect 4950 -4240 5550 -4120
rect 4950 -4480 5550 -4360
rect 4950 -4720 5550 -4600
rect 4950 -4960 5550 -4840
rect 4950 -5200 5550 -5080
rect 4950 -5440 5550 -5320
rect 4950 -5690 5550 -5560
rect 4950 -5930 5550 -5800
rect 4950 -6170 5550 -6050
<< nsubdiff >>
rect 4950 -900 5550 -870
rect 4950 -980 4980 -900
rect 5520 -980 5550 -900
rect 4950 -1000 5550 -980
rect 4670 -4540 4800 -4510
rect 4670 -5080 4690 -4540
rect 4770 -5080 4800 -4540
rect 4670 -5110 4800 -5080
<< nsubdiffcont >>
rect 4980 -980 5520 -900
rect 4690 -5080 4770 -4540
<< poly >>
rect 5690 -1020 5980 -1000
rect 5690 -1060 5710 -1020
rect 5750 -1040 5980 -1020
rect 5750 -1060 5770 -1040
rect 5690 -1080 5770 -1060
rect 4890 -1230 4950 -1110
rect 5550 -1230 5580 -1110
rect 4890 -1600 4920 -1230
rect 4890 -1720 4950 -1600
rect 5550 -1720 5580 -1600
rect 4890 -1840 4920 -1720
rect 4890 -1960 4950 -1840
rect 5550 -1960 5580 -1840
rect 4890 -2080 4920 -1960
rect 4890 -2200 4950 -2080
rect 5550 -2200 5580 -2080
rect 4890 -2320 4920 -2200
rect 4890 -2440 4950 -2320
rect 5550 -2440 5580 -2320
rect 5770 -2430 5850 -2410
rect 4890 -2560 4920 -2440
rect 5770 -2470 5790 -2430
rect 5830 -2450 5850 -2430
rect 5830 -2470 5990 -2450
rect 5770 -2490 5990 -2470
rect 4890 -2680 4950 -2560
rect 5550 -2680 5580 -2560
rect 4890 -2800 4920 -2680
rect 4890 -2920 4950 -2800
rect 5550 -2920 5580 -2800
rect 4890 -3040 4920 -2920
rect 4890 -3160 4950 -3040
rect 5550 -3160 5580 -3040
rect 4890 -3280 4920 -3160
rect 4890 -3400 4950 -3280
rect 5550 -3400 5580 -3280
rect 4890 -3760 4920 -3400
rect 4890 -3880 4950 -3760
rect 5550 -3880 5580 -3760
rect 4890 -4000 4920 -3880
rect 4890 -4120 4950 -4000
rect 5550 -4120 5580 -4000
rect 4890 -4240 4920 -4120
rect 4890 -4360 4950 -4240
rect 5550 -4360 5580 -4240
rect 4890 -4480 4920 -4360
rect 4890 -4600 4950 -4480
rect 5550 -4600 5580 -4480
rect 4890 -4720 4920 -4600
rect 4890 -4840 4950 -4720
rect 5550 -4840 5580 -4720
rect 4890 -4960 4920 -4840
rect 4890 -5080 4950 -4960
rect 5550 -5080 5580 -4960
rect 4890 -5200 4920 -5080
rect 4890 -5320 4950 -5200
rect 5550 -5320 5580 -5200
rect 4890 -5440 4920 -5320
rect 4890 -5560 4950 -5440
rect 5550 -5560 5580 -5440
rect 4890 -5930 4920 -5560
rect 4860 -6050 4950 -5930
rect 5550 -6050 5580 -5930
rect 4860 -6240 4890 -6050
rect 4860 -6260 4940 -6240
rect 4860 -6300 4880 -6260
rect 4920 -6300 4940 -6260
rect 4860 -6320 4940 -6300
<< polycont >>
rect 5710 -1060 5750 -1020
rect 5790 -2470 5830 -2430
rect 4880 -6300 4920 -6260
<< locali >>
rect 1820 -1160 2360 -1060
rect 1690 -1300 2410 -1220
rect 4060 -1950 4100 150
rect 5590 -850 5820 -830
rect 4960 -900 5540 -880
rect 4960 -980 4980 -900
rect 5520 -980 5540 -900
rect 4960 -1020 5540 -980
rect 4960 -1080 4980 -1020
rect 5520 -1080 5540 -1020
rect 4960 -1100 5540 -1080
rect 5590 -900 5620 -850
rect 5800 -900 5820 -850
rect 5590 -920 5820 -900
rect 5590 -990 5650 -920
rect 4960 -1260 5540 -1250
rect 4960 -1340 4980 -1260
rect 5520 -1340 5540 -1260
rect 4960 -1350 5540 -1340
rect 4870 -1590 5540 -1480
rect 4870 -1950 4910 -1590
rect 5590 -1730 5630 -990
rect 4960 -1830 5630 -1730
rect 2610 -1970 4910 -1950
rect 2610 -1990 5540 -1970
rect 2810 -2160 2920 -2060
rect 4870 -2070 5540 -1990
rect 4870 -2450 4910 -2070
rect 5590 -2210 5630 -1830
rect 4960 -2310 5630 -2210
rect 4870 -2550 5540 -2450
rect 4870 -2930 4910 -2550
rect 5590 -2690 5630 -2310
rect 4960 -2790 5630 -2690
rect 4870 -3030 5540 -2930
rect 4870 -3410 4910 -3030
rect 5590 -3170 5630 -2790
rect 4960 -3270 5630 -3170
rect 5690 -1020 5770 -1000
rect 5690 -1060 5710 -1020
rect 5750 -1060 5770 -1020
rect 5690 -1080 5770 -1060
rect 5690 -3310 5730 -1080
rect 5590 -3350 5730 -3310
rect 5770 -2430 5850 -2410
rect 5770 -2470 5790 -2430
rect 5830 -2470 5850 -2430
rect 5770 -2490 5850 -2470
rect 4870 -3510 5540 -3410
rect 4870 -3750 5540 -3650
rect 4870 -4130 4910 -3750
rect 5590 -3890 5630 -3350
rect 4960 -3990 5630 -3890
rect 4870 -4230 5540 -4130
rect 4670 -4540 4790 -4520
rect 2020 -5090 3930 -5050
rect 2020 -5200 2460 -5090
rect 3890 -6060 3930 -5090
rect 4670 -5080 4690 -4540
rect 4770 -5080 4790 -4540
rect 4670 -5100 4790 -5080
rect 4870 -4610 4910 -4230
rect 5590 -4370 5630 -3990
rect 4960 -4390 5630 -4370
rect 4960 -4450 4980 -4390
rect 5520 -4450 5630 -4390
rect 4960 -4470 5630 -4450
rect 4870 -4710 5540 -4610
rect 4870 -5090 4910 -4710
rect 5590 -4850 5630 -4470
rect 4960 -4950 5630 -4850
rect 4870 -5190 5540 -5090
rect 4870 -5570 4910 -5190
rect 5590 -5330 5630 -4950
rect 4960 -5430 5630 -5330
rect 4870 -5590 5540 -5570
rect 4870 -5660 4970 -5590
rect 5510 -5660 5540 -5590
rect 4870 -5670 5540 -5660
rect 4960 -5680 5540 -5670
rect 4960 -5830 5540 -5810
rect 4960 -5900 4980 -5830
rect 5520 -5900 5540 -5830
rect 4960 -5920 5540 -5900
rect 5770 -6060 5820 -2490
rect 3890 -6160 5820 -6060
rect 4860 -6260 4940 -6240
rect 4860 -6300 4880 -6260
rect 4920 -6280 4940 -6260
rect 11840 -6280 11880 -5050
rect 4920 -6300 11880 -6280
rect 4860 -6320 11880 -6300
<< viali >>
rect 4980 -980 5520 -900
rect 4980 -1080 5520 -1020
rect 5620 -900 5800 -850
rect 4980 -1340 5520 -1260
rect 2570 -1990 2610 -1950
rect 4690 -5080 4770 -4540
rect 4980 -4450 5520 -4390
rect 4970 -5660 5510 -5590
rect 4980 -5900 5520 -5830
<< metal1 >>
rect 4000 -860 4160 150
rect 1470 -1020 4160 -860
rect 5590 -840 5820 -830
rect 1470 -1350 1620 -1020
rect 4000 -1250 4160 -1020
rect 4950 -900 5550 -870
rect 4950 -980 4980 -900
rect 5520 -980 5550 -900
rect 4950 -990 5550 -980
rect 5590 -900 5620 -840
rect 5800 -900 5820 -840
rect 5590 -920 5820 -900
rect 5590 -990 5660 -920
rect 4950 -1020 5660 -990
rect 4950 -1080 4980 -1020
rect 5520 -1080 5660 -1020
rect 4950 -1110 5660 -1080
rect 4000 -1260 5540 -1250
rect 4000 -1340 4980 -1260
rect 5520 -1340 5540 -1260
rect 4000 -1350 5540 -1340
rect 1470 -1490 2630 -1350
rect 1490 -1510 2630 -1490
rect 2550 -1950 2630 -1930
rect 2550 -1990 2570 -1950
rect 2610 -1990 2630 -1950
rect 2550 -2430 2630 -1990
rect 5880 -3680 6020 -3330
rect 4190 -3820 6020 -3680
rect 4960 -4390 5550 -4370
rect 4960 -4450 4980 -4390
rect 5520 -4450 5550 -4390
rect 4960 -4470 5550 -4450
rect 4670 -4540 4800 -4510
rect 4670 -5080 4690 -4540
rect 4770 -5080 4800 -4540
rect 4670 -5110 4800 -5080
rect 3719 -5210 5782 -5208
rect 3719 -5310 6720 -5210
rect 3719 -5311 5782 -5310
rect 3720 -5380 3820 -5311
rect 2970 -5480 3820 -5380
rect 4960 -5590 5540 -5570
rect 4960 -5660 4970 -5590
rect 5510 -5660 5540 -5590
rect 4960 -5680 5540 -5660
rect 4960 -5830 5540 -5810
rect 4960 -5900 4980 -5830
rect 5520 -5900 5540 -5830
rect 4960 -5920 5540 -5900
<< via1 >>
rect 4980 -980 5520 -900
rect 5620 -850 5800 -840
rect 5620 -900 5800 -850
rect 4980 -1080 5520 -1020
rect 4980 -4450 5520 -4390
rect 4690 -5080 4770 -4540
rect 4970 -5660 5510 -5590
rect 4980 -5900 5520 -5830
<< metal2 >>
rect 5590 -840 5820 -830
rect 4950 -900 5550 -870
rect 4950 -980 4980 -900
rect 5520 -980 5550 -900
rect 4950 -990 5550 -980
rect 5590 -900 5620 -840
rect 5800 -900 5820 -840
rect 5590 -920 5820 -900
rect 5590 -990 5660 -920
rect 4950 -1020 5660 -990
rect 4950 -1080 4980 -1020
rect 5520 -1080 5660 -1020
rect 4950 -1110 5660 -1080
rect 5620 -1230 5660 -1110
rect 5620 -1290 6140 -1230
rect 2460 -3980 2540 -3660
rect 2460 -4020 4190 -3980
rect 4150 -4350 4190 -4020
rect 4150 -4390 5550 -4350
rect 4960 -4450 4980 -4390
rect 5520 -4450 5550 -4390
rect 4960 -4470 5550 -4450
rect 4670 -4540 4800 -4510
rect 4670 -5080 4690 -4540
rect 4770 -5080 4800 -4540
rect 4670 -5110 4800 -5080
rect 4960 -5590 5540 -5570
rect 4960 -5660 4970 -5590
rect 5510 -5660 5540 -5590
rect 4960 -5810 5540 -5660
rect 4960 -5830 5670 -5810
rect 4960 -5900 4980 -5830
rect 5520 -5900 5670 -5830
rect 4960 -5910 5670 -5900
rect 4960 -5920 5540 -5910
rect 5610 -6210 5670 -5910
rect 6370 -6210 6470 -5720
rect 5610 -6260 6470 -6210
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620692581
transform 1 0 6478 0 1 -10866
box -510 4630 8890 10940
<< end >>
