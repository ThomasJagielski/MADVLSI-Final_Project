**.subckt bandgap_pnp_lvs
XR2 __UNCONNECTED_PIN__0 __UNCONNECTED_PIN__1 GND sky130_fd_pr__res_xhigh_po W=0.35 L=3.5 mult=1 m=1
**.ends
.GLOBAL GND
** flattened .save nodes
.end
