**.subckt counter_lvs
X43 Qn0 __UNCONNECTED_PIN__0 net2 net1 P C dff
X44 net2 Qn0 __UNCONNECTED_PIN__1 net3 C P dff
X45 net1 net3 VDD GND inverter
X46 Qn1 __UNCONNECTED_PIN__2 net4 net12 P C dff
X53 net4 Qn1 __UNCONNECTED_PIN__3 Q0 C P dff
X54 Q0 net12 VDD GND inverter
X55 Qn2 __UNCONNECTED_PIN__4 net5 net13 P C dff
X56 net5 Qn2 __UNCONNECTED_PIN__5 Q1 C P dff
X57 Qn3 __UNCONNECTED_PIN__6 net6 net14 P C dff
X58 net6 Qn3 __UNCONNECTED_PIN__7 Q2 C P dff
X61 Q1 net13 VDD GND inverter
X62 Q2 net14 VDD GND inverter
X64 net2 Q0 VDD GND inverter
X65 net4 Q1 VDD GND inverter
X66 net5 Q2 VDD GND inverter
X67 net6 Q3 VDD GND inverter
X4 Qn4 __UNCONNECTED_PIN__8 net7 net15 P C dff
X5 net7 Qn4 __UNCONNECTED_PIN__9 Q3 C P dff
X7 Q3 net15 VDD GND inverter
X8 net7 Q4 VDD GND inverter
X9 Qn5 __UNCONNECTED_PIN__10 net8 net16 P C dff
X10 net8 Qn5 __UNCONNECTED_PIN__11 Q4 C P dff
X11 Q4 net16 VDD GND inverter
X12 Qn6 __UNCONNECTED_PIN__12 net9 net17 P C dff
X13 net9 Qn6 __UNCONNECTED_PIN__13 Q5 C P dff
X14 Qn7 __UNCONNECTED_PIN__14 net10 net18 P C dff
X15 net10 Qn7 __UNCONNECTED_PIN__15 Q6 C P dff
X18 Q5 net17 VDD GND inverter
X19 Q6 net18 VDD GND inverter
X21 net8 Q5 VDD GND inverter
X22 net9 Q6 VDD GND inverter
X23 net10 Q7 VDD GND inverter
X16 Qn8 __UNCONNECTED_PIN__16 net11 net19 P C dff
X17 net11 Qn8 __UNCONNECTED_PIN__17 Q7 C P dff
X20 Q7 net19 VDD GND inverter
X24 net11 Q8 VDD GND inverter
**.ends

* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/dff.sym # of pins=6

.subckt dff  D Qn Q CLK Preset Clear
*.ipin D
*.iopin CLK
*.opin Qn
*.opin Q
*.ipin Preset
*.ipin Clear
X6 D CLK net4 VDD GND nand2
X7 net1 CLK net2 VDD GND nand2
X8 Q net3 Qn VDD GND nand2
X9 net5 Qn Q VDD GND nand2
X10 D net1 VDD GND inverter
X1 VDD Preset GND net5 net4 and2
X2 VDD net2 GND net3 Clear and2
.ends


* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/inverter.sym # of
*+ pins=4

.subckt inverter  A Y VP VN
*.ipin A
*.iopin VP
*.iopin VN
*.opin Y
XM1 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 Y A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/nand2.sym # of pins=5

.subckt nand2  A B Y VP VN
*.ipin A
*.opin Y
*.ipin B
*.iopin VP
*.iopin VP
*.iopin VN
*.iopin VN
XM1 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 VP B Y VP sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net1 B Y VN sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net1 A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  /home/madvlsi/Documents/MADVLSI-Final_Project/schematic/and2.sym # of pins=5

.subckt and2  VP A VN Y B
*.iopin VP
*.iopin VN
*.ipin A
*.ipin B
*.opin Y
X1 A B net1 VP VN nand2
X2 net1 Y VP VN inverter
.ends

.GLOBAL VDD
.GLOBAL GND
** flattened .save nodes
.end
