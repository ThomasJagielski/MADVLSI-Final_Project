magic
tech sky130A
timestamp 1620776171
<< poly >>
rect 8780 1505 8825 1515
rect 8780 1485 8790 1505
rect 8815 1485 8825 1505
rect 8780 1475 8825 1485
rect 8785 -1760 8830 -1750
rect 8785 -1780 8795 -1760
rect 8820 -1780 8830 -1760
rect 8785 -1790 8830 -1780
rect 17615 -2560 17695 -2545
rect 17615 -2580 17625 -2560
rect 17645 -2580 17695 -2560
rect 17615 -2590 17695 -2580
<< polycont >>
rect 8790 1485 8815 1505
rect 8795 -1780 8820 -1760
rect 17625 -2580 17645 -2560
<< locali >>
rect 8780 1505 8825 1515
rect 8780 1485 8790 1505
rect 8815 1485 8825 1505
rect 8780 1475 8825 1485
rect 8980 1285 9085 1305
rect 8980 1215 9000 1285
rect 9065 1215 9085 1285
rect 8980 1180 9085 1215
rect 7345 1140 9085 1180
rect 7440 1100 7480 1110
rect 7290 1080 7450 1100
rect 7470 1080 7480 1100
rect 7290 1060 7480 1080
rect 8980 -385 9085 1140
rect 8980 -405 9260 -385
rect 17550 -1310 17610 -1300
rect 17550 -1325 17560 -1310
rect 15870 -1350 17560 -1325
rect 17600 -1350 17610 -1310
rect 17550 -1360 17610 -1350
rect 8600 -1435 9180 -1425
rect 8600 -1455 8610 -1435
rect 8630 -1455 9150 -1435
rect 9170 -1455 9180 -1435
rect 8600 -1465 9180 -1455
rect 8785 -1760 8830 -1750
rect 8785 -1780 8795 -1760
rect 8820 -1780 8830 -1760
rect 8785 -1790 8830 -1780
rect 17615 -2560 17655 -2545
rect 17615 -2580 17625 -2560
rect 17645 -2580 17655 -2560
rect 17615 -2590 17655 -2580
rect 17615 -2765 17695 -2755
rect 17615 -2795 17625 -2765
rect 17665 -2795 17695 -2765
rect 17615 -2805 17695 -2795
rect 8985 -3920 9090 -3900
rect 8985 -3990 9005 -3920
rect 9070 -3990 9090 -3920
rect 8985 -4300 9090 -3990
rect 7365 -4340 9090 -4300
<< viali >>
rect 8790 1485 8815 1505
rect 9000 1215 9065 1285
rect 7450 1080 7470 1100
rect 17560 -1350 17600 -1310
rect 8610 -1455 8630 -1435
rect 9150 -1455 9170 -1435
rect 8795 -1780 8820 -1760
rect 17625 -2580 17645 -2560
rect 17625 -2795 17665 -2765
rect 9005 -3990 9070 -3920
<< metal1 >>
rect 4610 5375 17695 5560
rect 4610 3305 4710 5375
rect 4610 3250 5620 3305
rect 4610 3075 4710 3250
rect 5520 3075 5620 3250
rect 8780 1510 8830 1515
rect 8780 1480 8785 1510
rect 8820 1480 8830 1510
rect 8780 1455 8830 1480
rect 7440 1435 8830 1455
rect 7440 1110 7460 1435
rect 7440 1100 7480 1110
rect 7240 1070 7290 1090
rect 7440 1080 7450 1100
rect 7470 1080 7480 1100
rect 7440 1070 7480 1080
rect 7365 -1425 7385 25
rect 8780 -100 8830 1435
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 13560 1060 13660 5375
rect 13560 865 13570 1060
rect 13650 865 13660 1060
rect 13560 580 13660 865
rect 8780 -135 10025 -100
rect 7365 -1435 8640 -1425
rect 7365 -1445 8610 -1435
rect 8600 -1455 8610 -1445
rect 8630 -1455 8640 -1435
rect 8600 -1465 8640 -1455
rect 8780 -1755 8830 -135
rect 17550 -1310 17610 -1300
rect 17550 -1350 17560 -1310
rect 17600 -1350 17610 -1310
rect 17550 -1360 17610 -1350
rect 9140 -1435 12755 -1425
rect 9140 -1455 9150 -1435
rect 9170 -1445 12755 -1435
rect 9170 -1455 9180 -1445
rect 9140 -1465 9180 -1455
rect 8780 -1785 8790 -1755
rect 8825 -1785 8830 -1755
rect 8780 -1790 8830 -1785
rect 8785 -1885 8830 -1825
rect 12720 -2120 12755 -1445
rect 12720 -2160 17655 -2120
rect 17615 -2560 17655 -2160
rect 17615 -2580 17625 -2560
rect 17645 -2580 17655 -2560
rect 17615 -2590 17655 -2580
rect 17615 -2765 17675 -2755
rect 17615 -2795 17625 -2765
rect 17665 -2795 17675 -2765
rect 17615 -2805 17675 -2795
rect 8995 -3920 9080 -3910
rect 8995 -3990 9005 -3920
rect 9070 -3990 9080 -3920
rect 8995 -4000 9080 -3990
rect 7405 -5485 18080 -5465
<< via1 >>
rect 8785 1505 8820 1510
rect 8785 1485 8790 1505
rect 8790 1485 8815 1505
rect 8815 1485 8820 1505
rect 8785 1480 8820 1485
rect 9000 1215 9065 1285
rect 13570 865 13650 1060
rect 17560 -1350 17600 -1310
rect 8790 -1760 8825 -1755
rect 8790 -1780 8795 -1760
rect 8795 -1780 8820 -1760
rect 8820 -1780 8825 -1760
rect 8790 -1785 8825 -1780
rect 17625 -2795 17665 -2765
rect 9005 -3990 9070 -3920
<< metal2 >>
rect 4005 5355 17695 5560
rect 4005 3075 4540 5355
rect 8780 1510 8825 1515
rect 8780 1480 8785 1510
rect 8820 1480 8825 1510
rect 8780 1475 8825 1480
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 12960 585 13395 5355
rect 13560 1060 13660 1070
rect 13560 865 13570 1060
rect 13650 865 13660 1060
rect 13560 855 13660 865
rect 7365 -1425 7385 25
rect 17550 -1310 17610 -1300
rect 17550 -1350 17560 -1310
rect 17600 -1350 17610 -1310
rect 17550 -1360 17610 -1350
rect 7365 -1445 12755 -1425
rect 8785 -1755 8830 -1750
rect 8785 -1785 8790 -1755
rect 8825 -1785 8830 -1755
rect 8785 -1790 8830 -1785
rect 12720 -2120 12755 -1445
rect 12720 -2160 17655 -2120
rect 17615 -2755 17655 -2160
rect 17615 -2765 17675 -2755
rect 17615 -2795 17625 -2765
rect 17665 -2795 17675 -2765
rect 17615 -2805 17675 -2795
rect 8995 -3920 9080 -3910
rect 8995 -3990 9005 -3920
rect 9070 -3990 9080 -3920
rect 8995 -4000 9080 -3990
rect 7405 -5485 18080 -5465
<< via2 >>
rect 8785 1480 8820 1510
rect 9000 1215 9065 1285
rect 13570 865 13650 1060
rect 17560 -1350 17600 -1310
rect 8790 -1785 8825 -1755
rect 9005 -3990 9070 -3920
<< metal3 >>
rect 8775 1510 8830 1585
rect 8775 1480 8785 1510
rect 8820 1480 8830 1510
rect 8775 1475 8830 1480
rect 8990 1285 9075 1295
rect 8990 1215 9000 1285
rect 9065 1215 9075 1285
rect 8990 1205 9075 1215
rect 12445 1060 13660 1070
rect 12445 865 13570 1060
rect 13650 865 13660 1060
rect 12445 855 13660 865
rect 17550 -1310 17695 -1300
rect 17550 -1350 17560 -1310
rect 17600 -1350 17695 -1310
rect 17550 -1360 17695 -1350
rect 8780 -1755 8835 -1750
rect 8780 -1785 8790 -1755
rect 8825 -1785 8835 -1755
rect 8780 -1855 8835 -1785
rect 8995 -3920 9080 -3910
rect 8995 -3990 9005 -3920
rect 9070 -3990 9080 -3920
rect 8995 -4000 9080 -3990
<< via3 >>
rect 9000 1215 9065 1285
rect 9005 -3990 9070 -3920
<< metal4 >>
rect 8980 1285 9085 1840
rect 8980 1215 9000 1285
rect 9065 1215 9085 1285
rect 8980 -1580 9085 1215
rect 8985 -2125 9090 -1580
rect 8985 -3920 9090 -3320
rect 8985 -3990 9005 -3920
rect 9070 -3990 9090 -3920
rect 8985 -4065 9090 -3990
use middle_ping_pong_amplifier  middle_ping_pong_amplifier_0
timestamp 1620710927
transform 1 0 12905 0 1 -1890
box -3700 -30 4680 3175
use bandgap_ping_pong_half  bandgap_ping_pong_half_0
timestamp 1620776171
transform 1 0 0 0 1 0
box -255 -5485 8650 5305
use cap8to1  cap8to1_1
timestamp 1620776171
transform 1 0 8760 0 1 1495
box 5 30 3785 1860
use cap8to1  cap8to1_0
timestamp 1620776171
transform 1 0 8765 0 1 -3670
box 5 30 3785 1860
<< end >>
