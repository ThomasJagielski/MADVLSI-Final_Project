magic
tech sky130A
timestamp 1620711011
<< nwell >>
rect -3180 2480 -2825 2725
rect -3175 1845 -2820 2090
<< nmos >>
rect -3110 2210 -3095 2310
rect -3035 2210 -3020 2410
rect -2960 2210 -2945 2310
rect -3105 1575 -3090 1675
rect -3030 1575 -3015 1775
rect -2955 1575 -2940 1675
<< pmos >>
rect -3110 2605 -3095 2705
rect -3035 2505 -3020 2705
rect -2960 2605 -2945 2705
rect -3105 1970 -3090 2070
rect -3030 1870 -3015 2070
rect -2955 1970 -2940 2070
<< ndiff >>
rect -3085 2395 -3035 2410
rect -3085 2310 -3070 2395
rect -3160 2295 -3110 2310
rect -3160 2225 -3145 2295
rect -3125 2225 -3110 2295
rect -3160 2210 -3110 2225
rect -3095 2225 -3070 2310
rect -3050 2225 -3035 2395
rect -3095 2210 -3035 2225
rect -3020 2395 -2970 2410
rect -3020 2225 -3005 2395
rect -2985 2310 -2970 2395
rect -2985 2225 -2960 2310
rect -3020 2210 -2960 2225
rect -2945 2295 -2895 2310
rect -2945 2225 -2930 2295
rect -2910 2225 -2895 2295
rect -2945 2210 -2895 2225
rect -3080 1760 -3030 1775
rect -3080 1675 -3065 1760
rect -3155 1660 -3105 1675
rect -3155 1590 -3140 1660
rect -3120 1590 -3105 1660
rect -3155 1575 -3105 1590
rect -3090 1590 -3065 1675
rect -3045 1590 -3030 1760
rect -3090 1575 -3030 1590
rect -3015 1760 -2965 1775
rect -3015 1590 -3000 1760
rect -2980 1675 -2965 1760
rect -2980 1590 -2955 1675
rect -3015 1575 -2955 1590
rect -2940 1660 -2890 1675
rect -2940 1590 -2925 1660
rect -2905 1590 -2890 1660
rect -2940 1575 -2890 1590
<< pdiff >>
rect -3160 2690 -3110 2705
rect -3160 2620 -3145 2690
rect -3125 2620 -3110 2690
rect -3160 2605 -3110 2620
rect -3095 2690 -3035 2705
rect -3095 2605 -3070 2690
rect -3085 2520 -3070 2605
rect -3050 2520 -3035 2690
rect -3085 2505 -3035 2520
rect -3020 2690 -2960 2705
rect -3020 2520 -3005 2690
rect -2985 2605 -2960 2690
rect -2945 2690 -2895 2705
rect -2945 2620 -2930 2690
rect -2910 2620 -2895 2690
rect -2945 2605 -2895 2620
rect -2985 2520 -2970 2605
rect -3020 2505 -2970 2520
rect -3155 2055 -3105 2070
rect -3155 1985 -3140 2055
rect -3120 1985 -3105 2055
rect -3155 1970 -3105 1985
rect -3090 2055 -3030 2070
rect -3090 1970 -3065 2055
rect -3080 1885 -3065 1970
rect -3045 1885 -3030 2055
rect -3080 1870 -3030 1885
rect -3015 2055 -2955 2070
rect -3015 1885 -3000 2055
rect -2980 1970 -2955 2055
rect -2940 2055 -2890 2070
rect -2940 1985 -2925 2055
rect -2905 1985 -2890 2055
rect -2940 1970 -2890 1985
rect -2980 1885 -2965 1970
rect -3015 1870 -2965 1885
<< ndiffc >>
rect -3145 2225 -3125 2295
rect -3070 2225 -3050 2395
rect -3005 2225 -2985 2395
rect -2930 2225 -2910 2295
rect -3140 1590 -3120 1660
rect -3065 1590 -3045 1760
rect -3000 1590 -2980 1760
rect -2925 1590 -2905 1660
<< pdiffc >>
rect -3145 2620 -3125 2690
rect -3070 2520 -3050 2690
rect -3005 2520 -2985 2690
rect -2930 2620 -2910 2690
rect -3140 1985 -3120 2055
rect -3065 1885 -3045 2055
rect -3000 1885 -2980 2055
rect -2925 1985 -2905 2055
<< psubdiff >>
rect -2935 2385 -2875 2400
rect -2935 2365 -2920 2385
rect -2890 2365 -2875 2385
rect -2935 2350 -2875 2365
rect -2930 1750 -2870 1765
rect -2930 1730 -2915 1750
rect -2885 1730 -2870 1750
rect -2930 1715 -2870 1730
<< nsubdiff >>
rect -2935 2540 -2875 2555
rect -2935 2520 -2920 2540
rect -2890 2520 -2875 2540
rect -2935 2505 -2875 2520
rect -2930 1905 -2870 1920
rect -2930 1885 -2915 1905
rect -2885 1885 -2870 1905
rect -2930 1870 -2870 1885
<< psubdiffcont >>
rect -2920 2365 -2890 2385
rect -2915 1730 -2885 1750
<< nsubdiffcont >>
rect -2920 2520 -2890 2540
rect -2915 1885 -2885 1905
<< poly >>
rect -3160 2750 -2945 2760
rect -3160 2730 -3150 2750
rect -3130 2745 -2945 2750
rect -3130 2730 -3095 2745
rect -3160 2720 -3095 2730
rect -3110 2705 -3095 2720
rect -3035 2705 -3020 2720
rect -2960 2705 -2945 2745
rect -2795 2735 -2750 2745
rect -2795 2715 -2785 2735
rect -2760 2715 -2750 2735
rect -2795 2705 -2750 2715
rect -1690 2710 -1645 2720
rect -3110 2590 -3095 2605
rect -1690 2690 -1680 2710
rect -1655 2690 -1645 2710
rect -1690 2680 -1645 2690
rect -3035 2490 -3020 2505
rect -3110 2475 -3020 2490
rect -3110 2310 -3095 2475
rect -2960 2465 -2945 2605
rect -100 2600 20 2615
rect -3000 2450 -2945 2465
rect -3000 2440 -2985 2450
rect -3035 2425 -2985 2440
rect -3035 2410 -3020 2425
rect -2960 2310 -2945 2425
rect -3110 2195 -3095 2210
rect -3035 2195 -3020 2210
rect -3160 2185 -3095 2195
rect -3160 2165 -3150 2185
rect -3130 2170 -3095 2185
rect -2960 2170 -2945 2210
rect -3130 2165 -2945 2170
rect -3160 2155 -2945 2165
rect -3155 2115 -2940 2125
rect -3155 2095 -3145 2115
rect -3125 2110 -2940 2115
rect -3125 2095 -3090 2110
rect -3155 2085 -3090 2095
rect -3105 2070 -3090 2085
rect -3030 2070 -3015 2085
rect -2955 2070 -2940 2110
rect -3105 1955 -3090 1970
rect -3030 1855 -3015 1870
rect -3105 1840 -3015 1855
rect -3105 1675 -3090 1840
rect -2955 1830 -2940 1970
rect -2995 1815 -2940 1830
rect -2995 1805 -2980 1815
rect -3030 1790 -2980 1805
rect -3030 1775 -3015 1790
rect -2955 1675 -2940 1790
rect -3105 1560 -3090 1575
rect -3030 1560 -3015 1575
rect -3155 1550 -3090 1560
rect -3155 1530 -3145 1550
rect -3125 1535 -3090 1550
rect -2955 1535 -2940 1575
rect -3125 1530 -2940 1535
rect -3155 1520 -2940 1530
rect -3525 1510 -3480 1520
rect -3525 1490 -3515 1510
rect -3490 1490 -3480 1510
rect -3525 1480 -3480 1490
rect -100 -335 -85 2600
rect -60 1880 5 1890
rect -60 1860 -50 1880
rect -30 1875 5 1880
rect -30 1860 -20 1875
rect -60 1850 -20 1860
rect -10 -335 35 -325
rect -100 -350 0 -335
rect -10 -355 0 -350
rect 25 -355 35 -335
rect -10 -365 35 -355
<< polycont >>
rect -3150 2730 -3130 2750
rect -2785 2715 -2760 2735
rect -1680 2690 -1655 2710
rect -3150 2165 -3130 2185
rect -3145 2095 -3125 2115
rect -3145 1530 -3125 1550
rect -3515 1490 -3490 1510
rect -50 1860 -30 1880
rect 0 -355 25 -335
<< locali >>
rect -2250 2785 -2145 2805
rect -3160 2750 -3120 2760
rect -3160 2730 -3150 2750
rect -3130 2730 -3120 2750
rect -3160 2720 -3120 2730
rect -2795 2735 -2750 2745
rect -2795 2715 -2785 2735
rect -2760 2715 -2750 2735
rect -3155 2690 -3040 2700
rect -3155 2620 -3145 2690
rect -3125 2620 -3070 2690
rect -3155 2610 -3070 2620
rect -3080 2520 -3070 2610
rect -3050 2520 -3040 2690
rect -3080 2475 -3040 2520
rect -3555 2425 -3480 2465
rect -3180 2435 -3040 2475
rect -3525 1830 -3480 2425
rect -3080 2395 -3040 2435
rect -3080 2305 -3070 2395
rect -3155 2295 -3070 2305
rect -3155 2225 -3145 2295
rect -3125 2225 -3070 2295
rect -3050 2225 -3040 2395
rect -3155 2215 -3040 2225
rect -3015 2690 -2895 2700
rect -3015 2520 -3005 2690
rect -2985 2620 -2930 2690
rect -2910 2620 -2895 2690
rect -2985 2610 -2895 2620
rect -2985 2520 -2975 2610
rect -3015 2475 -2975 2520
rect -2930 2540 -2880 2550
rect -2930 2520 -2920 2540
rect -2890 2520 -2880 2540
rect -2930 2510 -2880 2520
rect -2795 2475 -2750 2715
rect -2250 2715 -2230 2785
rect -2165 2715 -2145 2785
rect -2250 2695 -2145 2715
rect -1690 2710 -1645 2720
rect -3015 2435 -2750 2475
rect -3015 2395 -2975 2435
rect -3015 2225 -3005 2395
rect -2985 2305 -2975 2395
rect -2930 2385 -2880 2395
rect -2930 2365 -2920 2385
rect -2890 2365 -2880 2385
rect -2930 2355 -2880 2365
rect -2985 2295 -2895 2305
rect -2985 2225 -2930 2295
rect -2910 2225 -2895 2295
rect -3015 2215 -2895 2225
rect -3160 2185 -3120 2195
rect -3160 2165 -3150 2185
rect -3130 2165 -3120 2185
rect -3160 2155 -3120 2165
rect -3155 2115 -3115 2125
rect -3155 2095 -3145 2115
rect -3125 2095 -3115 2115
rect -3155 2085 -3115 2095
rect -3150 2055 -3035 2065
rect -3150 1985 -3140 2055
rect -3120 1985 -3065 2055
rect -3150 1975 -3065 1985
rect -3075 1885 -3065 1975
rect -3045 1885 -3035 2055
rect -3075 1840 -3035 1885
rect -3550 1790 -3480 1830
rect -3175 1800 -3035 1840
rect -3525 1510 -3480 1790
rect -3075 1760 -3035 1800
rect -3075 1670 -3065 1760
rect -3150 1660 -3065 1670
rect -3150 1590 -3140 1660
rect -3120 1590 -3065 1660
rect -3045 1590 -3035 1760
rect -3150 1580 -3035 1590
rect -3010 2055 -2890 2065
rect -3010 1885 -3000 2055
rect -2980 1985 -2925 2055
rect -2905 1985 -2890 2055
rect -2980 1975 -2890 1985
rect -2980 1885 -2970 1975
rect -3010 1840 -2970 1885
rect -2925 1905 -2875 1915
rect -2925 1885 -2915 1905
rect -2885 1885 -2875 1905
rect -2925 1875 -2875 1885
rect -2795 1840 -2750 2435
rect -3010 1800 -2750 1840
rect -2220 1890 -2175 2695
rect -1690 2690 -1680 2710
rect -1655 2690 -1645 2710
rect -1690 2680 -1645 2690
rect -2220 1880 -20 1890
rect -2220 1865 -50 1880
rect -2220 1830 -2175 1865
rect -60 1860 -50 1865
rect -30 1860 -20 1880
rect -60 1850 -20 1860
rect -3010 1760 -2970 1800
rect -2245 1790 -2175 1830
rect -3010 1590 -3000 1760
rect -2980 1670 -2970 1760
rect -2925 1750 -2875 1760
rect -2925 1730 -2915 1750
rect -2885 1730 -2875 1750
rect -2925 1720 -2875 1730
rect -2980 1660 -2890 1670
rect -2980 1590 -2925 1660
rect -2905 1590 -2890 1660
rect -3010 1580 -2890 1590
rect -3155 1550 -3115 1560
rect -3155 1530 -3145 1550
rect -3125 1530 -3115 1550
rect -3155 1520 -3115 1530
rect -3525 1490 -3515 1510
rect -3490 1490 -3480 1510
rect -3525 1480 -3480 1490
rect 2920 595 3130 610
rect 2875 570 3130 595
rect 2875 -45 2920 570
rect 725 -65 2920 -45
rect -10 -335 35 -325
rect -10 -355 0 -335
rect 25 -355 35 -335
rect -10 -415 35 -355
rect 685 -415 725 -395
rect -10 -445 725 -415
rect 2875 -425 2920 -65
rect 2815 -445 2920 -425
rect 2815 -515 2835 -445
rect 2900 -515 2920 -445
rect 2815 -535 2920 -515
<< viali >>
rect -2785 2715 -2760 2735
rect -2230 2715 -2165 2785
rect -1680 2690 -1655 2710
rect -3515 1490 -3490 1510
rect 0 -355 25 -335
rect 2835 -515 2900 -445
<< metal1 >>
rect -2240 2785 -2155 2795
rect -2795 2740 -2750 2745
rect -2795 2710 -2790 2740
rect -2755 2710 -2750 2740
rect -2795 2705 -2750 2710
rect -2240 2715 -2230 2785
rect -2165 2715 -2155 2785
rect -2240 2705 -2155 2715
rect -1690 2715 -1645 2720
rect -1690 2685 -1685 2715
rect -1650 2685 -1645 2715
rect -1690 2680 -1645 2685
rect -3525 1515 -3480 1520
rect -3525 1485 -3520 1515
rect -3485 1485 -3480 1515
rect -3525 1480 -3480 1485
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -10 -365 35 -360
rect 2825 -445 2910 -435
rect 2825 -515 2835 -445
rect 2900 -515 2910 -445
rect 2825 -525 2910 -515
<< via1 >>
rect -2790 2735 -2755 2740
rect -2790 2715 -2785 2735
rect -2785 2715 -2760 2735
rect -2760 2715 -2755 2735
rect -2790 2710 -2755 2715
rect -2230 2715 -2165 2785
rect -1685 2710 -1650 2715
rect -1685 2690 -1680 2710
rect -1680 2690 -1655 2710
rect -1655 2690 -1650 2710
rect -1685 2685 -1650 2690
rect -3520 1510 -3485 1515
rect -3520 1490 -3515 1510
rect -3515 1490 -3490 1510
rect -3490 1490 -3485 1510
rect -3520 1485 -3485 1490
rect -5 -335 30 -330
rect -5 -355 0 -335
rect 0 -355 25 -335
rect 25 -355 30 -335
rect -5 -360 30 -355
rect 2835 -515 2900 -445
<< metal2 >>
rect -2240 2785 -2155 2795
rect -2795 2740 -2750 2745
rect -2795 2710 -2790 2740
rect -2755 2710 -2750 2740
rect -2795 2705 -2750 2710
rect -2240 2715 -2230 2785
rect -2165 2715 -2155 2785
rect -2240 2705 -2155 2715
rect -1690 2715 -1645 2720
rect -1690 2685 -1685 2715
rect -1650 2685 -1645 2715
rect -1690 2680 -1645 2685
rect -3525 1515 -3480 1520
rect -3525 1485 -3520 1515
rect -3485 1485 -3480 1515
rect -3525 1480 -3480 1485
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -10 -365 35 -360
rect 2825 -445 2910 -435
rect 2825 -515 2835 -445
rect 2900 -515 2910 -445
rect 2825 -525 2910 -515
<< via2 >>
rect -2790 2710 -2755 2740
rect -2230 2715 -2165 2785
rect -1685 2685 -1650 2715
rect -3520 1485 -3485 1515
rect -5 -360 30 -330
rect 2835 -515 2900 -445
<< metal3 >>
rect -3020 3120 -2145 3220
rect -2800 2740 -2745 3025
rect -2800 2710 -2790 2740
rect -2755 2710 -2745 2740
rect -2800 2705 -2745 2710
rect -2240 2785 -2155 2795
rect -2240 2715 -2230 2785
rect -2165 2715 -2155 2785
rect -2240 2705 -2155 2715
rect -1695 2715 -1640 2975
rect -1695 2685 -1685 2715
rect -1650 2685 -1640 2715
rect -1695 2680 -1640 2685
rect -3525 1520 -3480 1570
rect -3530 1515 -3475 1520
rect -3530 1485 -3520 1515
rect -3485 1485 -3475 1515
rect -3530 1320 -3475 1485
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -1525 -520 -1430 -390
rect -10 -520 35 -360
rect -1525 -555 35 -520
rect 2825 -445 2910 -435
rect 2825 -515 2835 -445
rect 2900 -515 2910 -445
rect 2825 -525 2910 -515
<< via3 >>
rect -2230 2715 -2165 2785
rect 2835 -515 2900 -445
<< metal4 >>
rect -3020 3120 -2145 3220
rect -2250 2785 -2145 3120
rect -2250 2715 -2230 2785
rect -2165 2715 -2145 2785
rect -2250 2695 -2145 2715
rect -1755 -185 -985 -70
rect -1755 -425 -1630 -185
rect -1755 -445 2920 -425
rect -1755 -515 2835 -445
rect 2900 -515 2920 -445
rect -1755 -535 2920 -515
use switch  switch_4
timestamp 1620697026
transform 1 0 -2490 0 1 1490
box -110 20 245 625
use cap8to1  cap8to1_1
timestamp 1620709858
transform 1 0 -3890 0 1 2875
box 5 30 3785 1860
use switch  switch_3
timestamp 1620697026
transform 1 0 -3800 0 1 2125
box -110 20 245 625
use switch  switch_2
timestamp 1620697026
transform 1 0 -3795 0 1 1490
box -110 20 245 625
use switch  switch_1
timestamp 1620697026
transform 1 0 3170 0 1 270
box -110 20 245 625
use cap8to1  cap8to1_0
timestamp 1620709858
transform 1 0 -3915 0 1 -430
box 5 30 3785 1860
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620692581
transform 1 0 255 0 1 -2315
box -255 2315 4445 5470
use switch  switch_0
timestamp 1620697026
transform 0 -1 1025 1 0 -290
box -110 20 245 625
<< labels >>
rlabel locali -3160 2175 -3160 2175 7 nCLK
rlabel locali -3160 2740 -3160 2740 7 CLK
rlabel locali -2825 2455 -2825 2455 3 B
rlabel locali -3180 2455 -3180 2455 7 A
rlabel locali -3155 1540 -3155 1540 7 nCLK
rlabel locali -3155 2105 -3155 2105 7 CLK
rlabel locali -2820 1820 -2820 1820 3 B
rlabel locali -3175 1820 -3175 1820 7 A
rlabel locali -2245 1810 -2245 1810 3 B
<< end >>
