magic
tech sky130A
timestamp 1620435178
<< locali >>
rect 785 85 810 105
rect 0 65 120 85
rect 225 65 390 85
rect 495 65 660 85
rect 0 0 160 20
rect 430 -20 450 0
rect 0 -40 450 -20
use nand2  nand2_2
timestamp 1620350317
transform 1 0 660 0 1 60
box -120 -60 150 535
use nand2  nand2_1
timestamp 1620350317
transform 1 0 390 0 1 60
box -120 -60 150 535
use nand2  nand2_0
timestamp 1620350317
transform 1 0 120 0 1 60
box -120 -60 150 535
<< end >>
