magic
tech sky130A
timestamp 1620743260
<< poly >>
rect -85 -2000 -35 -1985
rect -85 -2020 -70 -2000
rect -50 -2020 -35 -2000
rect -85 -2125 -35 -2020
rect -85 -2145 -70 -2125
rect -50 -2145 -35 -2125
rect -85 -2160 -35 -2145
<< polycont >>
rect -70 -2020 -50 -2000
rect -70 -2145 -50 -2125
<< locali >>
rect -165 3390 55 3425
rect -165 -2055 -135 3390
rect -75 3000 35 3040
rect -75 -1985 -45 3000
rect -85 -2000 -35 -1985
rect -85 -2020 -70 -2000
rect -50 -2020 -35 -2000
rect -85 -2035 -35 -2020
rect -165 -2090 65 -2055
rect -85 -2125 -35 -2110
rect -85 -2145 -70 -2125
rect -50 -2145 -35 -2125
rect -85 -2440 -35 -2145
rect -85 -2480 50 -2440
<< metal1 >>
rect -235 3285 35 3325
rect -235 -2785 -200 3285
rect 6220 205 6770 930
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 6220 110 6770 120
rect -120 -5 25 15
rect -120 -2155 -75 -5
rect 6220 -90 6770 -80
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -970 6770 -175
rect 5335 -1505 6770 -970
rect 5335 -1975 5645 -1505
rect -120 -2195 45 -2155
rect 4625 -2285 5645 -1975
rect 4625 -2405 4725 -2285
rect 5545 -2405 5645 -2285
rect -235 -2820 25 -2785
<< via1 >>
rect 6230 120 6760 205
rect 6230 -175 6760 -90
<< metal2 >>
rect -235 2720 15 2760
rect -235 -3350 -200 2720
rect 4005 685 4425 835
rect 4005 470 4270 685
rect 4005 405 4015 470
rect 4260 405 4270 470
rect 4005 395 4270 405
rect 6220 205 6770 215
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 6220 110 6770 120
rect -120 -5 25 15
rect -120 -2720 -75 -5
rect 4025 -65 4355 -55
rect 4025 -145 4035 -65
rect 4345 -145 4355 -65
rect 4025 -2405 4355 -145
rect 6220 -90 6770 -80
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -185 6770 -175
rect -120 -2760 30 -2720
rect -235 -3390 60 -3350
<< via2 >>
rect 4015 405 4260 470
rect 6230 120 6760 205
rect 4035 -145 4345 -65
rect 6230 -175 6760 -90
<< metal3 >>
rect -250 3155 1405 3210
rect -250 -2270 -190 3155
rect 4005 470 4270 480
rect 4005 405 4015 470
rect 4260 405 4270 470
rect 4005 395 4270 405
rect 4025 -55 4270 395
rect 6220 205 6770 215
rect 6220 120 6230 205
rect 6760 120 6770 205
rect 4025 -65 4355 -55
rect 4025 -145 4035 -65
rect 4345 -145 4355 -65
rect 4025 -155 4355 -145
rect 6220 -90 6770 120
rect 6220 -175 6230 -90
rect 6760 -175 6770 -90
rect 6220 -185 6770 -175
rect -255 -2320 1260 -2270
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_1 ~/Documents/MADVLSI-Final_Project/layout
timestamp 1620741313
transform 1 0 3950 0 1 -4910
box -3935 -575 4700 4735
use bandgap_ping_pong_amp_cell  bandgap_ping_pong_amp_cell_0
timestamp 1620741313
transform 1 0 3930 0 1 570
box -3935 -575 4700 4735
<< end >>
