magic
tech sky130A
timestamp 1620773905
<< nwell >>
rect -3910 2715 -3850 2720
rect -3130 2715 -3090 2720
rect -3665 2500 -3605 2550
rect -3665 1870 -3555 1920
rect -3150 1885 -3040 1920
rect -3020 1885 -2975 1920
rect -2955 1885 -2845 1920
rect -3150 1870 -2845 1885
rect -2355 1870 -2295 1920
rect 3310 645 3360 685
rect 610 -150 650 -100
<< pmos >>
rect -3005 1870 -2990 1920
<< pdiff >>
rect -3055 1885 -3040 1920
rect -3020 1885 -3005 1920
rect -3055 1870 -3005 1885
rect -2990 1885 -2975 1920
rect -2955 1885 -2940 1920
rect -2990 1870 -2940 1885
<< psubdiff >>
rect -3660 2380 -3610 2390
rect -3660 2360 -3650 2380
rect -3620 2360 -3610 2380
rect -3660 2350 -3610 2360
rect -2900 2380 -2850 2390
rect -2900 2360 -2890 2380
rect -2860 2360 -2850 2380
rect -2900 2350 -2850 2360
rect -3660 1750 -3610 1760
rect -3660 1730 -3650 1750
rect -3620 1730 -3610 1750
rect -3660 1720 -3610 1730
rect -2900 1750 -2850 1760
rect -2900 1730 -2890 1750
rect -2860 1730 -2850 1750
rect -2900 1720 -2850 1730
<< nsubdiff >>
rect -3665 2535 -3605 2550
rect -3665 2515 -3650 2535
rect -3620 2515 -3605 2535
rect -3665 2500 -3605 2515
rect -3665 1905 -3605 1920
rect -3665 1885 -3650 1905
rect -3620 1885 -3605 1905
rect -3665 1870 -3605 1885
rect -2905 1905 -2845 1920
rect -2905 1885 -2890 1905
rect -2860 1885 -2845 1905
rect -2905 1870 -2845 1885
rect -2355 1905 -2295 1920
rect -2355 1885 -2340 1905
rect -2310 1885 -2295 1905
rect -2355 1870 -2295 1885
rect 3310 675 3360 685
rect 3310 655 3320 675
rect 3350 655 3360 675
rect 3310 645 3360 655
rect 610 -110 650 -100
rect 610 -140 620 -110
rect 640 -140 650 -110
rect 610 -150 650 -140
<< psubdiffcont >>
rect -3650 2360 -3620 2380
rect -2890 2360 -2860 2380
rect -3650 1730 -3620 1750
rect -2890 1730 -2860 1750
<< nsubdiffcont >>
rect -3650 2515 -3620 2535
rect -3650 1885 -3620 1905
rect -2890 1885 -2860 1905
rect -2340 1885 -2310 1905
rect 3320 655 3350 675
rect 620 -140 640 -110
<< poly >>
rect -2795 2905 -2750 2915
rect -2795 2885 -2785 2905
rect -2760 2885 -2750 2905
rect -2795 2875 -2750 2885
rect -3890 2745 -3850 2755
rect -3890 2725 -3880 2745
rect -3860 2725 -3850 2745
rect -3890 2715 -3850 2725
rect -3130 2745 -3090 2755
rect -3130 2725 -3120 2745
rect -3100 2725 -3090 2745
rect -3130 2715 -3090 2725
rect -1690 2710 -1645 2720
rect -1690 2690 -1680 2710
rect -1655 2690 -1645 2710
rect -1690 2680 -1645 2690
rect -100 2600 20 2615
rect -2630 2510 -2585 2520
rect -2630 2490 -2620 2510
rect -2600 2490 -2585 2510
rect -2630 2480 -2585 2490
rect -2630 2260 -2585 2270
rect -2630 2240 -2620 2260
rect -2600 2240 -2585 2260
rect -2630 2230 -2585 2240
rect -3890 2180 -3850 2190
rect -3890 2160 -3880 2180
rect -3860 2160 -3850 2180
rect -3890 2150 -3850 2160
rect -3130 2180 -3090 2190
rect -3130 2160 -3120 2180
rect -3100 2160 -3090 2180
rect -3130 2150 -3090 2160
rect -2930 1870 -2915 1920
rect -3130 1550 -3090 1560
rect -3130 1530 -3120 1550
rect -3100 1530 -3090 1550
rect -3130 1520 -3090 1530
rect -2580 1550 -2535 1560
rect -2580 1530 -2570 1550
rect -2550 1530 -2535 1550
rect -2580 1520 -2535 1530
rect -3525 1470 -3480 1480
rect -3525 1450 -3515 1470
rect -3490 1450 -3480 1470
rect -3525 1440 -3480 1450
rect -100 -520 -85 2600
rect -60 1880 5 1890
rect -60 1860 -50 1880
rect -30 1875 5 1880
rect -30 1860 -20 1875
rect -60 1850 -20 1860
rect 620 -445 725 -425
rect 620 -515 640 -445
rect 705 -515 725 -445
rect 620 -520 725 -515
rect -100 -535 725 -520
<< polycont >>
rect -2785 2885 -2760 2905
rect -3880 2725 -3860 2745
rect -3120 2725 -3100 2745
rect -1680 2690 -1655 2710
rect -2620 2490 -2600 2510
rect -2620 2240 -2600 2260
rect -3880 2160 -3860 2180
rect -3120 2160 -3100 2180
rect -3120 2095 -3100 2115
rect -3120 1530 -3100 1550
rect -2570 1530 -2550 1550
rect -3515 1450 -3490 1470
rect -50 1860 -30 1880
rect 975 -370 995 -350
rect 640 -515 705 -445
<< locali >>
rect -2795 2905 -2750 2915
rect -2795 2885 -2785 2905
rect -2760 2885 -2750 2905
rect -3915 2820 -3275 2855
rect -3890 2745 -3850 2755
rect -3890 2725 -3880 2745
rect -3860 2725 -3850 2745
rect -3890 2715 -3850 2725
rect -3660 2540 -3610 2545
rect -3660 2510 -3650 2540
rect -3620 2510 -3610 2540
rect -3660 2505 -3610 2510
rect -3310 2470 -3275 2820
rect -3130 2745 -3090 2755
rect -3130 2725 -3120 2745
rect -3100 2725 -3090 2745
rect -3130 2715 -3090 2725
rect -2795 2475 -2750 2885
rect -2250 2785 -2145 2805
rect -2250 2715 -2230 2785
rect -2165 2715 -2145 2785
rect -2250 2695 -2145 2715
rect -1690 2710 -1645 2720
rect -2630 2510 -2590 2520
rect -2630 2490 -2620 2510
rect -2600 2490 -2590 2510
rect -2630 2480 -2590 2490
rect -3555 2430 -3480 2470
rect -3310 2430 -3140 2470
rect -2800 2435 -2750 2475
rect -3660 2380 -3610 2390
rect -3660 2360 -3650 2380
rect -3620 2360 -3610 2380
rect -3660 2350 -3610 2360
rect -3890 2180 -3850 2190
rect -3890 2160 -3880 2180
rect -3860 2160 -3850 2180
rect -3890 2150 -3850 2160
rect -3660 1910 -3610 1915
rect -3660 1880 -3650 1910
rect -3620 1880 -3610 1910
rect -3660 1875 -3610 1880
rect -3525 1840 -3480 2430
rect -2900 2380 -2850 2390
rect -2900 2360 -2890 2380
rect -2860 2360 -2850 2380
rect -2900 2350 -2850 2360
rect -3130 2180 -3090 2190
rect -3130 2160 -3120 2180
rect -3100 2160 -3090 2180
rect -3130 2150 -3090 2160
rect -3050 1885 -3040 1920
rect -3020 1885 -3010 1920
rect -3050 1870 -3010 1885
rect -2985 1885 -2975 1920
rect -2955 1885 -2945 1920
rect -2985 1870 -2945 1885
rect -2900 1910 -2850 1915
rect -2900 1880 -2890 1910
rect -2860 1880 -2850 1910
rect -2900 1875 -2850 1880
rect -2795 1840 -2750 2435
rect -2630 2260 -2590 2270
rect -2630 2240 -2620 2260
rect -2600 2240 -2590 2260
rect -2630 2230 -2590 2240
rect -2350 1910 -2300 1915
rect -2350 1880 -2340 1910
rect -2310 1880 -2300 1910
rect -2350 1875 -2300 1880
rect -2220 1890 -2175 2695
rect -1690 2690 -1680 2710
rect -1655 2690 -1645 2710
rect -1690 2680 -1645 2690
rect -2220 1880 -20 1890
rect -2220 1865 -50 1880
rect -2220 1840 -2175 1865
rect -60 1860 -50 1865
rect -30 1860 -20 1880
rect -60 1850 -20 1860
rect -3935 1800 -3885 1840
rect -3555 1800 -3480 1840
rect -3935 1415 -3910 1800
rect -3660 1750 -3610 1760
rect -3660 1730 -3650 1750
rect -3620 1730 -3610 1750
rect -3660 1720 -3610 1730
rect -3525 1470 -3480 1800
rect -3235 1825 -3145 1840
rect -3235 1805 -3220 1825
rect -3200 1805 -3145 1825
rect -3235 1800 -3145 1805
rect -2800 1800 -2750 1840
rect -2685 1800 -2570 1840
rect -2245 1800 -2175 1840
rect -3235 1790 -3165 1800
rect -3525 1450 -3515 1470
rect -3490 1450 -3480 1470
rect -3525 1440 -3480 1450
rect -3185 1495 -3165 1790
rect -2900 1750 -2850 1760
rect -2900 1730 -2890 1750
rect -2860 1730 -2850 1750
rect -2900 1720 -2850 1730
rect -3130 1550 -3090 1560
rect -3130 1530 -3120 1550
rect -3100 1530 -3090 1550
rect -3130 1520 -3090 1530
rect -2685 1495 -2660 1800
rect -2580 1550 -2540 1560
rect -2580 1530 -2570 1550
rect -2550 1530 -2540 1550
rect -2580 1520 -2540 1530
rect -3185 1465 -2660 1495
rect -3185 1415 -3165 1465
rect -3935 1395 -3165 1415
rect 3080 885 3120 895
rect 3080 865 3090 885
rect 3110 865 3120 885
rect 3080 855 3120 865
rect 3310 680 3360 685
rect 3310 650 3320 680
rect 3350 650 3360 680
rect 3310 645 3360 650
rect 2875 570 3130 610
rect 2875 -25 2920 570
rect -10 -50 2920 -25
rect -10 -335 35 -50
rect 610 -110 650 -100
rect 610 -140 615 -110
rect 645 -140 650 -110
rect 610 -150 650 -140
rect -10 -355 0 -335
rect 25 -355 35 -335
rect 965 -350 1005 -340
rect -10 -365 35 -355
rect 965 -370 975 -350
rect 995 -370 1005 -350
rect 965 -380 1005 -370
rect 685 -425 725 -390
rect 620 -445 725 -425
rect 620 -515 640 -445
rect 705 -515 725 -445
rect 620 -535 725 -515
<< viali >>
rect -2785 2885 -2760 2905
rect -3880 2725 -3860 2745
rect -3650 2535 -3620 2540
rect -3650 2515 -3620 2535
rect -3650 2510 -3620 2515
rect -3120 2725 -3100 2745
rect -2890 2510 -2860 2540
rect -2230 2715 -2165 2785
rect -2620 2490 -2600 2510
rect -3650 2360 -3620 2380
rect -3880 2160 -3860 2180
rect -3880 2095 -3860 2115
rect -3650 1905 -3620 1910
rect -3650 1885 -3620 1905
rect -3650 1880 -3620 1885
rect -2890 2360 -2860 2380
rect -3120 2160 -3100 2180
rect -3120 2095 -3100 2115
rect -2890 1905 -2860 1910
rect -2890 1885 -2860 1905
rect -2890 1880 -2860 1885
rect -2620 2240 -2600 2260
rect -2570 2095 -2550 2115
rect -2340 1905 -2310 1910
rect -2340 1885 -2310 1905
rect -2340 1880 -2310 1885
rect -1680 2690 -1655 2710
rect -3650 1730 -3620 1750
rect -3880 1530 -3860 1550
rect -3220 1805 -3200 1825
rect -3515 1450 -3490 1470
rect -2890 1730 -2860 1750
rect -3120 1530 -3100 1550
rect -2340 1730 -2310 1750
rect -2570 1530 -2550 1550
rect 3090 865 3110 885
rect 3320 675 3350 680
rect 3320 655 3350 675
rect 3320 650 3350 655
rect 3320 500 3350 520
rect 3090 300 3110 320
rect 615 -140 620 -110
rect 620 -140 640 -110
rect 640 -140 645 -110
rect 775 -140 795 -110
rect 0 -355 25 -335
rect 410 -370 430 -350
rect 975 -370 995 -350
rect 640 -515 705 -445
<< metal1 >>
rect -2795 2910 -2750 2915
rect -2795 2880 -2790 2910
rect -2755 2880 -2750 2910
rect -2795 2875 -2750 2880
rect -2240 2785 -2155 2795
rect -3910 2745 -2600 2755
rect -3910 2725 -3880 2745
rect -3860 2725 -3120 2745
rect -3100 2725 -2600 2745
rect -3910 2715 -2600 2725
rect -3660 2540 -3610 2545
rect -3660 2510 -3650 2540
rect -3620 2510 -3610 2540
rect -3660 2505 -3610 2510
rect -2900 2540 -2850 2545
rect -2900 2510 -2890 2540
rect -2860 2510 -2850 2540
rect -2620 2520 -2600 2715
rect -2240 2715 -2230 2785
rect -2165 2715 -2155 2785
rect -2240 2705 -2155 2715
rect -1690 2715 -1645 2720
rect -1690 2685 -1685 2715
rect -1650 2685 -1645 2715
rect -1690 2680 -1645 2685
rect -2900 2505 -2850 2510
rect -2630 2515 -2590 2520
rect -2630 2485 -2625 2515
rect -2595 2485 -2590 2515
rect -2630 2480 -2590 2485
rect -3660 2380 -3610 2390
rect -2900 2380 -2850 2390
rect -3660 2360 -3650 2380
rect -3620 2360 -2890 2380
rect -2860 2360 -2155 2380
rect -3660 2350 -3610 2360
rect -2900 2350 -2850 2360
rect -3890 2185 -3850 2190
rect -3890 2155 -3885 2185
rect -3855 2155 -3850 2185
rect -3890 2150 -3850 2155
rect -3130 2185 -3090 2190
rect -3130 2155 -3125 2185
rect -3095 2155 -3090 2185
rect -3130 2150 -3090 2155
rect -3930 2115 -3090 2125
rect -3930 2095 -3880 2115
rect -3860 2095 -3120 2115
rect -3100 2095 -3090 2115
rect -3930 2085 -3090 2095
rect -3930 -555 -3910 2085
rect -3660 1910 -3610 1915
rect -3660 1880 -3650 1910
rect -3620 1880 -3610 1910
rect -3660 1875 -3610 1880
rect -2900 1910 -2850 1915
rect -2900 1880 -2890 1910
rect -2860 1880 -2850 1910
rect -2900 1875 -2850 1880
rect -3235 1830 -3185 1840
rect -3235 1800 -3225 1830
rect -3195 1800 -3185 1830
rect -3235 1790 -3185 1800
rect -3660 1750 -3610 1760
rect -2900 1750 -2850 1760
rect -2750 1750 -2730 2360
rect -2620 2270 -2600 2275
rect -2630 2265 -2590 2270
rect -2630 2235 -2625 2265
rect -2595 2235 -2590 2265
rect -2630 2230 -2590 2235
rect -3660 1730 -3650 1750
rect -3620 1730 -2890 1750
rect -2860 1730 -2730 1750
rect -2620 2115 -2600 2230
rect -2580 2115 -2540 2125
rect -2620 2095 -2570 2115
rect -2550 2095 -2540 2115
rect -3660 1720 -3610 1730
rect -2900 1720 -2850 1730
rect -3890 1555 -3850 1560
rect -3890 1525 -3885 1555
rect -3855 1525 -3850 1555
rect -3890 1520 -3850 1525
rect -3130 1555 -3090 1560
rect -3130 1525 -3125 1555
rect -3095 1525 -3090 1555
rect -3130 1520 -3090 1525
rect -2620 1485 -2600 2095
rect -2580 2085 -2540 2095
rect -2175 2065 -2155 2360
rect -2175 2045 120 2065
rect -2350 1910 -2300 1915
rect -2350 1880 -2340 1910
rect -2310 1880 -2300 1910
rect -2350 1875 -2300 1880
rect -2350 1750 -2300 1760
rect -2175 1750 -2155 2045
rect -2350 1730 -2340 1750
rect -2310 1730 -2155 1750
rect -2350 1720 -2300 1730
rect -2580 1555 -2540 1560
rect -2580 1525 -2575 1555
rect -2545 1525 -2540 1555
rect -2580 1520 -2540 1525
rect -3525 1475 -3480 1480
rect -3525 1445 -3520 1475
rect -3485 1445 -3480 1475
rect -2620 1465 -95 1485
rect -3525 1440 -3480 1445
rect -115 -285 -95 1465
rect 3080 885 3120 895
rect 3080 865 3090 885
rect 3110 865 3455 885
rect 3080 855 3120 865
rect 3310 680 3360 685
rect 3310 650 3320 680
rect 3350 650 3360 680
rect 3310 645 3360 650
rect 3310 520 3360 530
rect 2790 500 3320 520
rect 3350 500 3360 520
rect 3310 490 3360 500
rect 3080 325 3120 330
rect 3080 295 3085 325
rect 3115 295 3120 325
rect 3080 290 3120 295
rect 690 -25 720 175
rect 690 -45 795 -25
rect 775 -100 795 -45
rect 610 -110 650 -100
rect 610 -140 615 -110
rect 645 -140 650 -110
rect 610 -150 650 -140
rect 765 -110 805 -100
rect 765 -140 775 -110
rect 795 -140 805 -110
rect 765 -150 805 -140
rect -115 -305 75 -285
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -10 -365 35 -360
rect 55 -405 75 -305
rect 400 -350 440 -340
rect 400 -370 410 -350
rect 430 -370 440 -350
rect 400 -405 440 -370
rect 965 -345 1005 -340
rect 965 -375 970 -345
rect 1000 -375 1005 -345
rect 965 -380 1005 -375
rect 55 -425 440 -405
rect 630 -445 715 -435
rect 630 -515 640 -445
rect 705 -515 715 -445
rect 630 -525 715 -515
rect 3435 -555 3455 865
rect -3930 -575 3455 -555
<< via1 >>
rect -2790 2905 -2755 2910
rect -2790 2885 -2785 2905
rect -2785 2885 -2760 2905
rect -2760 2885 -2755 2905
rect -2790 2880 -2755 2885
rect -3650 2510 -3620 2540
rect -2890 2510 -2860 2540
rect -2230 2715 -2165 2785
rect -1685 2710 -1650 2715
rect -1685 2690 -1680 2710
rect -1680 2690 -1655 2710
rect -1655 2690 -1650 2710
rect -1685 2685 -1650 2690
rect -2625 2510 -2595 2515
rect -2625 2490 -2620 2510
rect -2620 2490 -2600 2510
rect -2600 2490 -2595 2510
rect -2625 2485 -2595 2490
rect -3885 2180 -3855 2185
rect -3885 2160 -3880 2180
rect -3880 2160 -3860 2180
rect -3860 2160 -3855 2180
rect -3885 2155 -3855 2160
rect -3125 2180 -3095 2185
rect -3125 2160 -3120 2180
rect -3120 2160 -3100 2180
rect -3100 2160 -3095 2180
rect -3125 2155 -3095 2160
rect -3650 1880 -3620 1910
rect -2890 1880 -2860 1910
rect -3225 1825 -3195 1830
rect -3225 1805 -3220 1825
rect -3220 1805 -3200 1825
rect -3200 1805 -3195 1825
rect -3225 1800 -3195 1805
rect -2625 2260 -2595 2265
rect -2625 2240 -2620 2260
rect -2620 2240 -2600 2260
rect -2600 2240 -2595 2260
rect -2625 2235 -2595 2240
rect -3885 1550 -3855 1555
rect -3885 1530 -3880 1550
rect -3880 1530 -3860 1550
rect -3860 1530 -3855 1550
rect -3885 1525 -3855 1530
rect -3125 1550 -3095 1555
rect -3125 1530 -3120 1550
rect -3120 1530 -3100 1550
rect -3100 1530 -3095 1550
rect -3125 1525 -3095 1530
rect -2340 1880 -2310 1910
rect -2575 1550 -2545 1555
rect -2575 1530 -2570 1550
rect -2570 1530 -2550 1550
rect -2550 1530 -2545 1550
rect -2575 1525 -2545 1530
rect -3520 1470 -3485 1475
rect -3520 1450 -3515 1470
rect -3515 1450 -3490 1470
rect -3490 1450 -3485 1470
rect -3520 1445 -3485 1450
rect 3320 650 3350 680
rect 3085 320 3115 325
rect 3085 300 3090 320
rect 3090 300 3110 320
rect 3110 300 3115 320
rect 3085 295 3115 300
rect 615 -140 645 -110
rect -5 -335 30 -330
rect -5 -355 0 -335
rect 0 -355 25 -335
rect 25 -355 30 -335
rect -5 -360 30 -355
rect 970 -350 1000 -345
rect 970 -370 975 -350
rect 975 -370 995 -350
rect 995 -370 1000 -350
rect 970 -375 1000 -370
rect 640 -515 705 -445
<< metal2 >>
rect -2795 2910 -2750 2915
rect -2795 2880 -2790 2910
rect -2755 2880 -2750 2910
rect -2795 2875 -2750 2880
rect -2240 2785 -2155 2795
rect -2240 2715 -2230 2785
rect -2165 2715 -2155 2785
rect -2240 2705 -2155 2715
rect -1690 2715 -1645 2720
rect -1690 2685 -1685 2715
rect -1650 2685 -1645 2715
rect -1690 2680 -1645 2685
rect -3660 2540 -3610 2545
rect -3660 2535 -3650 2540
rect -3665 2515 -3650 2535
rect -3660 2510 -3650 2515
rect -3620 2535 -3610 2540
rect -2900 2540 -2850 2545
rect -2900 2535 -2890 2540
rect -3620 2515 -2890 2535
rect -3620 2510 -3610 2515
rect -3660 2505 -3610 2510
rect -2900 2510 -2890 2515
rect -2860 2535 -2850 2540
rect -2860 2515 -2660 2535
rect -2630 2520 -2585 2525
rect -2860 2510 -2850 2515
rect -2900 2505 -2850 2510
rect -2680 2385 -2660 2515
rect -2635 2480 -2630 2520
rect -2590 2480 -2585 2520
rect -2680 2365 130 2385
rect -3130 2190 -3085 2195
rect -3930 2185 -3130 2190
rect -3930 2155 -3885 2185
rect -3855 2155 -3130 2185
rect -3930 2150 -3130 2155
rect -3090 2150 -3085 2190
rect -3660 1910 -3610 1915
rect -3660 1905 -3650 1910
rect -3665 1885 -3650 1905
rect -3660 1880 -3650 1885
rect -3620 1905 -3610 1910
rect -2900 1910 -2850 1915
rect -2900 1905 -2890 1910
rect -3620 1885 -2890 1905
rect -3620 1880 -3610 1885
rect -3660 1875 -3610 1880
rect -2900 1880 -2890 1885
rect -2860 1905 -2850 1910
rect -2680 1905 -2660 2365
rect -2630 2270 -2585 2275
rect -2635 2230 -2630 2270
rect -2590 2230 -2585 2270
rect -2350 1910 -2300 1915
rect -2350 1905 -2340 1910
rect -2860 1885 -2340 1905
rect -2860 1880 -2850 1885
rect -2900 1875 -2850 1880
rect -2350 1880 -2340 1885
rect -2310 1905 -2300 1910
rect -2310 1885 -2295 1905
rect -2310 1880 -2300 1885
rect -2350 1875 -2300 1880
rect -3235 1830 -3185 1840
rect -3235 1800 -3225 1830
rect -3195 1800 -3185 1830
rect -3235 1790 -3185 1800
rect -2580 1560 -2535 1565
rect -3930 1555 -3090 1560
rect -3930 1525 -3885 1555
rect -3855 1525 -3125 1555
rect -3095 1525 -3090 1555
rect -3930 1520 -3090 1525
rect -2585 1520 -2580 1560
rect -2540 1550 -2535 1560
rect -2540 1530 -95 1550
rect -2540 1520 -2535 1530
rect -3930 -555 -3910 1520
rect -3525 1475 -3480 1480
rect -3525 1445 -3520 1475
rect -3485 1445 -3480 1475
rect -3525 1440 -3480 1445
rect -115 -285 -95 1530
rect 3310 680 3360 685
rect 3310 675 3320 680
rect 2990 655 3320 675
rect 450 -30 480 250
rect 2130 40 2160 140
rect 2990 40 3010 655
rect 3310 650 3320 655
rect 3350 650 3360 680
rect 3310 645 3360 650
rect 3080 325 3120 330
rect 3080 295 3085 325
rect 3115 320 3120 325
rect 3115 300 3455 320
rect 3115 295 3120 300
rect 3080 290 3120 295
rect 2130 20 3010 40
rect 450 -50 640 -30
rect 620 -100 640 -50
rect 610 -110 650 -100
rect 610 -140 615 -110
rect 645 -140 650 -110
rect 610 -150 650 -140
rect -115 -305 75 -285
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -10 -365 35 -360
rect 55 -350 75 -305
rect 965 -345 1005 -340
rect 965 -350 970 -345
rect 55 -370 970 -350
rect 965 -375 970 -370
rect 1000 -375 1005 -345
rect 965 -380 1005 -375
rect 630 -445 715 -435
rect 630 -515 640 -445
rect 705 -515 715 -445
rect 630 -525 715 -515
rect 3435 -555 3455 300
rect -3930 -575 3455 -555
<< via2 >>
rect -2790 2880 -2755 2910
rect -2230 2715 -2165 2785
rect -1685 2685 -1650 2715
rect -2630 2515 -2590 2520
rect -2630 2485 -2625 2515
rect -2625 2485 -2595 2515
rect -2595 2485 -2590 2515
rect -2630 2480 -2590 2485
rect -3130 2185 -3090 2190
rect -3130 2155 -3125 2185
rect -3125 2155 -3095 2185
rect -3095 2155 -3090 2185
rect -3130 2150 -3090 2155
rect -2630 2265 -2590 2270
rect -2630 2235 -2625 2265
rect -2625 2235 -2595 2265
rect -2595 2235 -2590 2265
rect -2630 2230 -2590 2235
rect -3225 1800 -3195 1830
rect -2580 1555 -2540 1560
rect -2580 1525 -2575 1555
rect -2575 1525 -2545 1555
rect -2545 1525 -2540 1555
rect -2580 1520 -2540 1525
rect -3520 1445 -3485 1475
rect -5 -360 30 -330
rect 640 -515 705 -445
<< metal3 >>
rect -3020 3120 -2715 3220
rect -2575 3120 -2145 3220
rect -2800 2910 -2745 3025
rect -2800 2880 -2790 2910
rect -2755 2880 -2745 2910
rect -2800 2875 -2745 2880
rect -2240 2785 -2155 2795
rect -2240 2715 -2230 2785
rect -2165 2715 -2155 2785
rect -2240 2705 -2155 2715
rect -1695 2715 -1640 2975
rect -1695 2685 -1685 2715
rect -1650 2685 -1640 2715
rect -1695 2640 -1640 2685
rect -3235 2590 -1640 2640
rect -3235 1830 -3185 2590
rect -2625 2525 -2595 2540
rect -2635 2520 -2585 2525
rect -2635 2480 -2630 2520
rect -2590 2480 -2585 2520
rect -2635 2475 -2585 2480
rect -2625 2275 -2595 2475
rect -2635 2270 -2585 2275
rect -2635 2230 -2630 2270
rect -2590 2230 -2585 2270
rect -2635 2225 -2585 2230
rect -3135 2190 -2190 2195
rect -3135 2150 -3130 2190
rect -3090 2150 -2190 2190
rect -3135 2145 -2190 2150
rect -3235 1800 -3225 1830
rect -3195 1800 -3185 1830
rect -3235 1790 -3185 1800
rect -3525 1480 -3480 1570
rect -2585 1560 -2535 1565
rect -2220 1560 -2190 2145
rect -2585 1520 -2580 1560
rect -2540 1520 -2190 1560
rect -2585 1515 -2535 1520
rect -3530 1475 -3475 1480
rect -3530 1445 -3520 1475
rect -3485 1445 -3475 1475
rect -3530 1320 -3475 1445
rect -10 -330 35 -325
rect -10 -360 -5 -330
rect 30 -360 35 -330
rect -1525 -520 -1430 -390
rect -10 -520 35 -360
rect -1525 -555 35 -520
rect 630 -445 715 -435
rect 630 -515 640 -445
rect 705 -515 715 -445
rect 630 -525 715 -515
<< via3 >>
rect -2230 2715 -2165 2785
rect 640 -515 705 -445
<< metal4 >>
rect -3020 3120 -2145 3220
rect -2250 2785 -2145 3120
rect -2250 2715 -2230 2785
rect -2165 2715 -2145 2785
rect -2250 2695 -2145 2715
rect -1755 -185 -985 -70
rect -1755 -425 -1630 -185
rect -1755 -445 725 -425
rect -1755 -515 640 -445
rect 705 -515 725 -445
rect -1755 -535 725 -515
use switch  switch_4
timestamp 1620697026
transform 1 0 -2490 0 1 1500
box -110 20 245 625
use switch  switch_2
timestamp 1620697026
transform 1 0 -3800 0 1 1500
box -110 20 245 625
use switch  switch_5
timestamp 1620697026
transform 1 0 -3040 0 1 1500
box -110 20 245 625
use switch  switch_3
timestamp 1620697026
transform 1 0 -3800 0 1 2130
box -110 20 245 625
use switch  switch_6
timestamp 1620697026
transform 1 0 -3040 0 1 2130
box -110 20 245 625
use switch  switch_0
timestamp 1620697026
transform 0 -1 1025 1 0 -290
box -110 20 245 625
use switch  switch_1
timestamp 1620697026
transform 1 0 3170 0 1 270
box -110 20 245 625
use cap8to1  cap8to1_0
timestamp 1620772218
transform 1 0 -3915 0 1 -430
box 5 30 3785 1860
use cap8to1  cap8to1_1
timestamp 1620772218
transform 1 0 -3890 0 1 2875
box 5 30 3785 1860
use selfbiasedcascode2stage  selfbiasedcascode2stage_0
timestamp 1620772218
transform 1 0 255 0 1 -2315
box -255 2315 4445 5470
<< labels >>
rlabel metal1 -3910 2735 -3910 2735 7 Vphi1
rlabel metal2 -3930 2170 -3930 2170 7 Vnphi1
rlabel metal1 -3930 2105 -3930 2105 7 Vphi2
rlabel metal1 -3930 1540 -3930 1540 7 Vnphi2
rlabel space -3910 2450 -3910 2450 7 Vn
rlabel locali -3915 2835 -3915 2835 7 Vp
<< end >>
